magic
tech sky130A
timestamp 1639202694
<< nwell >>
rect -16 301 140 519
<< nmos >>
rect 53 142 71 242
<< pmos >>
rect 53 360 71 460
<< ndiff >>
rect 3 229 53 242
rect 3 211 20 229
rect 37 211 53 229
rect 3 173 53 211
rect 3 155 20 173
rect 37 155 53 173
rect 3 142 53 155
rect 71 229 121 242
rect 71 211 87 229
rect 104 211 121 229
rect 71 173 121 211
rect 71 155 87 173
rect 104 155 121 173
rect 71 142 121 155
<< pdiff >>
rect 3 447 53 460
rect 3 429 20 447
rect 37 429 53 447
rect 3 391 53 429
rect 3 373 20 391
rect 37 373 53 391
rect 3 360 53 373
rect 71 447 121 460
rect 71 429 87 447
rect 104 429 121 447
rect 71 391 121 429
rect 71 373 87 391
rect 104 373 121 391
rect 71 360 121 373
<< ndiffc >>
rect 20 211 37 229
rect 20 155 37 173
rect 87 211 104 229
rect 87 155 104 173
<< pdiffc >>
rect 20 429 37 447
rect 20 373 37 391
rect 87 429 104 447
rect 87 373 104 391
<< poly >>
rect 45 502 79 510
rect 45 484 53 502
rect 71 484 79 502
rect 45 474 79 484
rect 53 460 71 474
rect 53 346 71 360
rect 45 336 79 346
rect 45 318 53 336
rect 71 318 79 336
rect 45 282 79 318
rect 45 264 53 282
rect 71 264 79 282
rect 45 256 79 264
rect 53 242 71 256
rect 53 128 71 142
rect 45 120 79 128
rect 45 102 53 120
rect 71 102 79 120
rect 45 94 79 102
<< polycont >>
rect 53 484 71 502
rect 53 318 71 336
rect 53 264 71 282
rect 53 102 71 120
<< locali >>
rect 45 509 79 510
rect 45 482 47 509
rect 77 482 79 509
rect 45 474 79 482
rect 10 450 46 456
rect 10 423 15 450
rect 10 420 46 423
rect 78 447 114 456
rect 78 429 87 447
rect 104 429 114 447
rect 78 420 114 429
rect 10 391 46 400
rect 10 373 20 391
rect 37 373 46 391
rect 10 364 46 373
rect 78 395 114 400
rect 78 368 83 395
rect 78 364 114 368
rect 45 336 79 346
rect 45 318 53 336
rect 71 318 79 336
rect 45 317 79 318
rect 45 290 47 317
rect 77 290 79 317
rect 45 282 79 290
rect 45 264 53 282
rect 71 264 79 282
rect 45 256 79 264
rect 10 229 46 238
rect 10 211 20 229
rect 37 211 46 229
rect 10 202 46 211
rect 78 229 114 238
rect 78 211 87 229
rect 104 211 114 229
rect 78 202 114 211
rect 10 178 46 182
rect 10 151 11 178
rect 42 151 46 178
rect 10 146 46 151
rect 78 178 114 182
rect 78 151 83 178
rect 78 146 114 151
rect 45 122 79 128
rect 45 95 47 122
rect 77 95 79 122
rect 45 94 79 95
<< viali >>
rect 47 502 77 509
rect 47 484 53 502
rect 53 484 71 502
rect 71 484 77 502
rect 47 482 77 484
rect 15 447 46 450
rect 15 429 20 447
rect 20 429 37 447
rect 37 429 46 447
rect 15 423 46 429
rect 83 391 114 395
rect 83 373 87 391
rect 87 373 104 391
rect 104 373 114 391
rect 83 368 114 373
rect 47 290 77 317
rect 11 173 42 178
rect 11 155 20 173
rect 20 155 37 173
rect 37 155 42 173
rect 11 151 42 155
rect 83 173 114 178
rect 83 155 87 173
rect 87 155 104 173
rect 104 155 114 173
rect 83 151 114 155
rect 47 120 77 122
rect 47 102 53 120
rect 53 102 71 120
rect 71 102 77 120
rect 47 95 77 102
<< metal1 >>
rect -328 465 -163 587
rect 41 509 84 514
rect 41 482 47 509
rect 77 482 84 509
rect 41 475 84 482
rect -328 454 -77 465
rect -6 454 51 459
rect -328 450 334 454
rect -328 426 15 450
rect -328 422 -77 426
rect -6 423 15 426
rect 46 426 334 450
rect 46 423 51 426
rect -328 -50 -163 422
rect -6 416 51 423
rect 78 395 135 402
rect 78 387 83 395
rect -89 368 83 387
rect 114 387 135 395
rect 114 368 335 387
rect -89 359 335 368
rect 41 317 84 322
rect 41 290 47 317
rect 77 290 84 317
rect 41 283 84 290
rect 1111 254 1130 298
rect -102 188 -30 195
rect -102 164 -98 188
rect -109 130 -98 164
rect -41 171 -30 188
rect -10 178 47 184
rect -10 171 11 178
rect -41 151 11 171
rect 42 151 47 178
rect -41 142 47 151
rect 77 178 134 185
rect 77 151 83 178
rect 114 170 134 178
rect 114 151 334 170
rect 77 142 334 151
rect -41 130 -30 142
rect -10 141 47 142
rect -109 123 -30 130
rect -109 119 -69 123
rect 41 122 84 127
rect 41 95 47 122
rect 77 95 84 122
rect 41 88 84 95
rect -328 -93 -77 -50
rect -328 -553 -163 -93
rect 1096 -253 1126 -214
rect -102 -330 -30 -323
rect -102 -388 -95 -330
rect -38 -388 -30 -330
rect -102 -395 -30 -388
rect -328 -596 -70 -553
rect -328 -1053 -163 -596
rect 1096 -762 1126 -723
rect -98 -833 -26 -826
rect -98 -891 -91 -833
rect -34 -891 -26 -833
rect -98 -898 -26 -891
rect -328 -1096 -77 -1053
rect -328 -1469 -163 -1096
rect 1096 -1265 1126 -1226
rect -98 -1329 -26 -1322
rect -98 -1387 -91 -1329
rect -34 -1387 -26 -1329
rect -98 -1394 -26 -1387
rect -266 -1489 -235 -1469
rect -266 -1520 274 -1489
rect -266 -1544 -235 -1520
rect -303 -1554 -235 -1544
rect 243 -1554 274 -1520
rect -303 -1585 -116 -1554
rect 243 -1585 357 -1554
rect -303 -1602 -248 -1585
rect -303 -1930 -272 -1602
rect 321 -1900 387 -1863
rect 321 -1915 813 -1900
rect 366 -1922 813 -1915
rect -303 -1961 350 -1930
rect -303 -2012 -272 -1961
rect -303 -2043 -113 -2012
rect 319 -2048 350 -1961
rect 369 -1970 813 -1922
rect 743 -2151 813 -1970
rect -142 -2180 -131 -2175
rect -149 -2189 -131 -2180
rect -149 -2199 -135 -2189
rect -143 -2239 -113 -2200
rect 612 -2221 813 -2151
rect 314 -2261 344 -2222
<< via1 >>
rect 47 482 77 509
rect 47 290 77 317
rect -98 130 -41 188
rect 47 95 77 122
rect -95 -388 -38 -330
rect -91 -891 -34 -833
rect -91 -1387 -34 -1329
rect -142 -1743 -111 -1707
rect 166 -1741 198 -1710
rect 336 -1736 376 -1706
rect 629 -1751 660 -1712
rect -123 -2192 -91 -2160
rect 181 -2204 210 -2176
rect 332 -2203 367 -2167
<< metal2 >>
rect 41 509 84 561
rect 41 482 47 509
rect 77 482 84 509
rect 41 475 84 482
rect 41 317 84 322
rect 41 290 47 317
rect 77 290 84 317
rect 41 283 84 290
rect -102 188 -30 198
rect -102 164 -98 188
rect -109 130 -98 164
rect -41 130 -30 188
rect -109 126 -30 130
rect -109 119 -69 126
rect 41 122 84 127
rect 41 95 47 122
rect 77 95 84 122
rect 41 48 84 95
rect 162 47 206 560
rect -105 -330 -33 -323
rect -105 -388 -95 -330
rect -38 -388 -33 -330
rect -105 -395 -33 -388
rect -98 -833 -26 -826
rect -98 -891 -91 -833
rect -34 -891 -26 -833
rect -98 -898 -26 -891
rect -98 -1329 -26 -1322
rect -98 -1387 -91 -1329
rect -34 -1387 -26 -1329
rect -98 -1394 -26 -1387
rect -162 -1471 84 -1427
rect -162 -1627 -118 -1471
rect -161 -1694 -118 -1627
rect -161 -1707 -100 -1694
rect 162 -1699 205 -1427
rect 331 -1470 503 -1427
rect 581 -1470 725 -1426
rect 331 -1690 374 -1470
rect 681 -1689 725 -1470
rect -161 -1736 -142 -1707
rect -150 -1743 -142 -1736
rect -111 -1743 -100 -1707
rect -150 -1750 -100 -1743
rect 154 -1710 210 -1699
rect 154 -1741 166 -1710
rect 198 -1741 210 -1710
rect 154 -1750 210 -1741
rect 320 -1706 394 -1690
rect 667 -1698 725 -1689
rect 320 -1736 336 -1706
rect 376 -1736 394 -1706
rect 320 -1748 394 -1736
rect 614 -1712 725 -1698
rect -150 -1754 -102 -1750
rect -150 -1898 -121 -1754
rect 324 -1765 359 -1748
rect 614 -1751 629 -1712
rect 660 -1751 725 -1712
rect 614 -1754 725 -1751
rect 614 -1764 672 -1754
rect -150 -1927 210 -1898
rect -143 -2151 -102 -2126
rect -143 -2160 -80 -2151
rect -143 -2172 -123 -2160
rect -133 -2192 -123 -2172
rect -91 -2192 -80 -2160
rect 181 -2162 210 -1927
rect 324 -2151 359 -2137
rect -133 -2201 -80 -2192
rect 172 -2176 224 -2162
rect 172 -2204 181 -2176
rect 210 -2204 224 -2176
rect 172 -2211 224 -2204
rect 320 -2167 391 -2151
rect 320 -2203 332 -2167
rect 367 -2203 391 -2167
rect 320 -2212 391 -2203
<< via2 >>
rect -98 130 -41 188
rect -95 -388 -38 -330
rect -91 -891 -34 -833
rect -91 -1387 -34 -1329
<< metal3 >>
rect -614 203 -371 602
rect -614 188 -27 203
rect -614 130 -98 188
rect -41 130 -27 188
rect -614 117 -27 130
rect -614 -317 -371 117
rect -614 -330 -20 -317
rect -614 -388 -95 -330
rect -38 -388 -20 -330
rect -614 -403 -20 -388
rect -614 -822 -371 -403
rect -614 -826 -27 -822
rect -614 -833 -26 -826
rect -614 -891 -91 -833
rect -34 -891 -26 -833
rect -614 -898 -26 -891
rect -614 -908 -27 -898
rect -614 -1320 -371 -908
rect -614 -1322 -27 -1320
rect -614 -1329 -26 -1322
rect -614 -1387 -91 -1329
rect -34 -1387 -26 -1329
rect -614 -1394 -26 -1387
rect -614 -1406 -27 -1394
rect -614 -1468 -371 -1406
rect 754 -1468 929 542
rect -623 -1516 929 -1468
rect -623 -1644 926 -1516
rect -131 -1820 -81 -1644
rect 247 -1818 297 -1644
rect -131 -1861 -73 -1820
rect -131 -1868 -90 -1861
rect 247 -1868 402 -1818
rect -123 -1914 -90 -1868
rect -123 -2200 -73 -1914
rect -143 -2239 -73 -2200
rect -123 -2326 -73 -2239
rect 336 -2332 386 -1868
use 0_unit  0_unit_2
timestamp 1639199462
transform 1 0 419 0 1 -1518
box -89 47 335 561
use 1  1_3
timestamp 1639199554
transform 1 0 0 0 1 -1518
box -89 47 335 561
use 1  1_2
timestamp 1639199554
transform 1 0 0 0 1 -1016
box -89 47 335 561
use 1  1_1
timestamp 1639199554
transform 1 0 420 0 1 -1016
box -89 47 335 561
use inv_customized  inv_customized_3
timestamp 1639194575
transform 1 0 933 0 1 -1520
box -194 128 180 481
use 0_unit  0_unit_1
timestamp 1639199462
transform 1 0 0 0 1 -512
box -89 47 335 561
use 1  1_0
timestamp 1639199554
transform 1 0 420 0 1 -512
box -89 47 335 561
use inv_customized  inv_customized_2
timestamp 1639194575
transform 1 0 933 0 1 -1018
box -194 128 180 481
use 0_unit  0_unit_0
timestamp 1639199462
transform 1 0 420 0 1 -1
box -89 47 335 561
use inv_customized  inv_customized_1
timestamp 1639194575
transform 1 0 937 0 1 -513
box -194 128 180 481
use inv_customized  inv_customized_0
timestamp 1639194575
transform 1 0 943 0 1 -1
box -194 128 180 481
use inv_customized  inv_customized_7
timestamp 1639194575
transform 1 0 502 0 1 -2474
box -194 128 180 481
use inv_customized  inv_customized_6
timestamp 1639194575
transform 1 0 47 0 1 -2468
box -194 128 180 481
use inv_customized  inv_customized_5
timestamp 1639194575
transform 1 0 35 0 1 -2010
box -194 128 180 481
use inv_customized  inv_customized_4
timestamp 1639194575
transform 1 0 498 0 1 -2010
box -194 128 180 481
<< labels >>
rlabel locali 62 290 62 290 5 Gate
port 1 n
rlabel viali 62 508 62 508 1 Gate
port 1 n
rlabel viali 62 313 62 313 1 Gate
port 2 n
rlabel metal2 60 560 60 560 1 N1
rlabel metal2 185 559 185 559 1 N2
rlabel metal1 -87 440 -87 440 7 W1
rlabel metal1 -88 371 -88 371 7 W2
rlabel via1 -88 156 -88 156 7 W3
rlabel metal1 333 440 333 440 3 E1
rlabel metal1 334 373 334 373 3 E2
rlabel metal1 333 157 333 157 3 E3
rlabel metal2 183 48 183 48 5 S2
rlabel metal2 61 49 61 49 5 S1
rlabel locali 63 95 63 95 1 Gate
port 2 s
rlabel metal3 -493 592 -493 592 1 GND
rlabel metal1 -248 570 -248 570 1 VDD
rlabel metal1 321 -2236 321 -2236 1 A0
rlabel metal1 1101 -1235 1101 -1235 1 sel3
rlabel metal1 1108 -738 1108 -738 1 sel2
rlabel metal1 1105 -236 1105 -236 1 sel1
rlabel metal1 1120 276 1120 276 7 sel0
rlabel metal1 -140 -2190 -140 -2190 1 A1
<< end >>
