* SPICE3 file created from 2x4_circuit.ext - technology: sky130A

.subckt x1 W3 S1 S2 SUB W1 W2 E3
X0 W1 S1 W2 w_106_301# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X1 W3 S1 E3 SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
.ends

.subckt inv_customized GND IN VDD SUB
X0 OUT IN VDD w_n16_301# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X1 OUT IN GND SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
.ends

.subckt x0_unit W3 S1 S2 SUB W1 W2 E3
X0 W2 S1 W1 w_n16_301# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X1 E3 S1 W3 SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
.ends

.subckt x2x4_circuit Gate
X1_0 1_0/W3 1_1/S1 1_1/S2 SUB W1 1_0/W3 1_0/E3 x1
X1_1 1_2/W2 1_1/S1 1_1/S2 SUB W1 1_2/W2 1_2/W3 x1
X1_2 1_2/W3 S2 Gate SUB W1 1_2/W2 W3 x1
X1_3 1_3/W3 S2 Gate SUB W1 1_3/W2 W3 x1
Xinv_customized_0 W3 W2 W1 SUB inv_customized
Xinv_customized_1 W3 1_0/W3 W1 SUB inv_customized
X0_unit_0 E3 1_1/S2 1_1/S1 SUB W1 W2 W2 x0_unit
Xinv_customized_2 W3 1_2/W2 W1 SUB inv_customized
X0_unit_1 W3 Gate S2 SUB W1 1_0/W3 1_0/E3 x0_unit
Xinv_customized_3 W3 1_3/W2 W1 SUB inv_customized
X0_unit_2 1_3/W3 1_1/S2 1_1/S1 SUB W1 1_3/W2 1_3/W2 x0_unit
X0 W2 Gate W1 w_n16_301# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X1 E3 Gate W3 SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
C0 W1 SUB -3.62fF
C1 W3 SUB -2.96fF
.ends

