* SPICE3 file created from 2x4_circuit.ext - technology: sky130A

.subckt x1 E1 E2 E3 W3 N1 N2 w_106_301# SUB
X0 E1 N1 E2 w_106_301# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X1 W3 N1 E3 SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
.ends

.subckt inv_customized VDD IN GND OUT SUB w_n16_301#
X0 OUT IN VDD w_n16_301# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X1 OUT IN GND SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
.ends

.subckt x0_unit W1 W2 W3 E3 N2 N1 SUB w_n16_301#
X0 W2 N1 W1 w_n16_301# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X1 E3 N1 W3 SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
.ends

.subckt x2x4_circuit Gate
X1_0 W1 1_0/W3 1_0/E3 1_0/W3 1_1/N1 1_1/N2 W1 W3 x1
X1_1 W1 1_2/E2 1_2/W3 1_2/E2 1_1/N1 1_1/N2 W1 W3 x1
X1_2 W1 1_2/E2 W3 1_2/W3 S2 Gate W1 W3 x1
X1_3 W1 1_3/E2 W3 1_3/W3 S2 Gate W1 W3 x1
Xinv_customized_0 W1 W2 W3 sel0 W3 W1 inv_customized
X0_unit_0 W1 W2 E3 W2 1_1/N1 1_1/N2 W3 W1 x0_unit
Xinv_customized_1 W1 1_0/W3 W3 sel1 W3 W1 inv_customized
X0_unit_1 W1 1_0/W3 W3 1_0/E3 S2 Gate W3 W1 x0_unit
Xinv_customized_2 W1 1_2/E2 W3 sel2 W3 W1 inv_customized
Xinv_customized_3 W1 1_3/E2 W3 sel3 W3 W1 inv_customized
X0_unit_2 W1 1_3/E2 1_3/W3 1_3/E2 1_1/N1 1_1/N2 W3 W1 x0_unit
Xinv_customized_4 W1 1_1/N2 W3 1_1/N1 W3 W1 inv_customized
Xinv_customized_5 W1 Gate W3 S2 W3 W1 inv_customized
Xinv_customized_6 W1 A1 W3 Gate W3 W1 inv_customized
Xinv_customized_7 W1 A0 W3 1_1/N2 W3 W1 inv_customized
X0 W2 Gate W1 W1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X1 E3 Gate W3 W3 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
C0 1_1/N2 W3 -3.24fF
C1 S2 W3 -2.37fF
C2 Gate W3 -4.38fF
C3 W1 W3 -16.74fF
C4 1_1/N1 W3 -2.77fF
.ends

