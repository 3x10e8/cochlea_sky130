magic
tech sky130A
timestamp 1639205400
use 0  0_23
timestamp 1639200303
transform -1 0 -178 0 1 -3658
box -89 43 336 566
use 0  0_22
timestamp 1639200303
transform -1 0 -178 0 1 -3135
box -89 43 336 566
use 0  0_18
timestamp 1639200303
transform 1 0 0 0 1 -3658
box -89 43 336 566
use 0  0_16
timestamp 1639200303
transform 1 0 0 0 1 -3135
box -89 43 336 566
use 0  0_19
timestamp 1639200303
transform 1 0 425 0 1 -3658
box -89 43 336 566
use 0  0_17
timestamp 1639200303
transform -1 0 672 0 1 -3135
box -89 43 336 566
use inv_customized  inv_customized_7
timestamp 1639201766
transform 1 0 951 0 1 -3661
box -194 128 180 481
use 0  0_21
timestamp 1639200303
transform -1 0 -178 0 1 -2612
box -89 43 336 566
use 0  0_15
timestamp 1639200303
transform -1 0 247 0 1 -2612
box -89 43 336 566
use 0  0_14
timestamp 1639200303
transform -1 0 672 0 1 -2612
box -89 43 336 566
use inv_customized  inv_customized_6
timestamp 1639201766
transform 1 0 951 0 1 -3138
box -194 128 180 481
use 0  0_20
timestamp 1639200303
transform -1 0 -178 0 1 -2089
box -89 43 336 566
use 0  0_12
timestamp 1639200303
transform -1 0 247 0 1 -2089
box -89 43 336 566
use 0  0_13
timestamp 1639200303
transform 1 0 425 0 1 -2089
box -89 43 336 566
use inv_customized  inv_customized_5
timestamp 1639201766
transform 1 0 951 0 1 -2615
box -194 128 180 481
use 0  0_11
timestamp 1639200303
transform 1 0 -425 0 1 -1566
box -89 43 336 566
use 0  0_2
timestamp 1639200303
transform -1 0 247 0 1 -1566
box -89 43 336 566
use 0  0_7
timestamp 1639200303
transform 1 0 425 0 1 -1566
box -89 43 336 566
use inv_customized  inv_customized_4
timestamp 1639201766
transform 1 0 951 0 1 -2092
box -194 128 180 481
use 0  0_10
timestamp 1639200303
transform 1 0 -425 0 1 -1043
box -89 43 336 566
use 0  0_4
timestamp 1639200303
transform -1 0 247 0 1 -1043
box -89 43 336 566
use 0  0_6
timestamp 1639200303
transform -1 0 672 0 1 -1043
box -89 43 336 566
use inv_customized  inv_customized_3
timestamp 1639201766
transform 1 0 951 0 1 -1569
box -194 128 180 481
use 0  0_9
timestamp 1639200303
transform 1 0 -425 0 1 -520
box -89 43 336 566
use 0  0_3
timestamp 1639200303
transform 1 0 0 0 1 -520
box -89 43 336 566
use 0  0_5
timestamp 1639200303
transform -1 0 672 0 1 -520
box -89 43 336 566
use inv_customized  inv_customized_2
timestamp 1639201766
transform 1 0 951 0 1 -1046
box -194 128 180 481
use 0  0_8
timestamp 1639200303
transform 1 0 -425 0 1 3
box -89 43 336 566
use 0  0_0
timestamp 1639200303
transform 1 0 0 0 1 3
box -89 43 336 566
use 0  0_1
timestamp 1639200303
transform 1 0 425 0 1 3
box -89 43 336 566
use inv_customized  inv_customized_1
timestamp 1639201766
transform 1 0 951 0 1 -523
box -194 128 180 481
use inv_customized  inv_customized_0
timestamp 1639201766
transform 1 0 951 0 1 0
box -194 128 180 481
<< end >>
