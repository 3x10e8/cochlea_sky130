* SPICE3 file created from 5x32.ext - technology: sky130A

.subckt x0 W1 W2 W3 E3 N2 N1 SUB w_n16_301#
X0 W2 N1 W1 w_n16_301# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X1 E3 N1 W3 SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
.ends

.subckt inv_customized VDD IN GND OUT SUB w_n16_301#
X0 OUT IN VDD w_n16_301# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X1 OUT IN GND SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
.ends

.subckt inv_customized_3 OUT GND IN VDD SUB w_n16_301#
X0 OUT IN VDD w_n16_301# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X1 OUT IN GND SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
.ends

.subckt x5x32 W1 W3
X0_138 W1 0_158/W2 0_139/E3 0_138/E3 0_9/N2 0_9/N1 W3 W1 x0
X0_127 W1 0_155/W2 0_155/W3 0_127/E3 0_97/N1 0_97/N2 W3 W1 x0
X0_116 W1 0_153/W2 0_153/W2 0_117/E3 0_7/N1 0_7/N2 W3 W1 x0
X0_105 W1 0_150/W2 0_106/W3 0_105/E3 0_4/N1 0_4/N2 W3 W1 x0
X0_149 W1 0_149/W2 0_149/W3 W3 0_79/N1 0_79/N2 W3 W1 x0
Xinv_customized_14 W1 0_72/W2 W3 inv_customized_14/OUT W3 W1 inv_customized
Xinv_customized_25 W1 0_151/W2 W3 inv_customized_25/OUT W3 W1 inv_customized
X0_139 W1 0_158/W2 0_158/W3 0_139/E3 0_97/N1 0_97/N2 W3 W1 x0
X0_128 W1 0_156/W2 0_131/W3 0_156/W2 0_7/N2 0_7/N1 W3 W1 x0
X0_117 W1 0_153/W2 0_118/W3 0_117/E3 0_4/N1 0_4/N2 W3 W1 x0
X0_106 W1 0_150/W2 0_106/W3 0_107/W3 0_9/N1 0_9/N2 W3 W1 x0
Xinv_customized_15 W1 0_79/W2 W3 inv_customized_15/OUT W3 W1 inv_customized
Xinv_customized_26 W1 0_99/W2 W3 inv_customized_26/OUT W3 W1 inv_customized
X0_129 W1 0_156/W2 0_130/E3 0_131/E3 0_9/N2 0_9/N1 W3 W1 x0
X0_118 W1 0_153/W2 0_118/W3 0_119/E3 0_9/N1 0_9/N2 W3 W1 x0
X0_107 W1 0_150/W2 0_107/W3 0_150/W3 0_97/N2 0_97/N1 W3 W1 x0
Xinv_customized_27 W1 0_149/W2 W3 inv_customized_27/OUT W3 W1 inv_customized
Xinv_customized_16 W1 0_159/W2 W3 inv_customized_16/OUT W3 W1 inv_customized
X0_119 W1 0_153/W2 0_153/W3 0_119/E3 0_97/N1 0_97/N2 W3 W1 x0
X0_108 W1 0_151/W2 0_109/E3 0_151/W2 0_7/N2 0_7/N1 W3 W1 x0
Xinv_customized_28 W1 0_91/W2 W3 inv_customized_28/OUT W3 W1 inv_customized
Xinv_customized_17 W1 0_158/W2 W3 inv_customized_17/OUT W3 W1 inv_customized
X0_109 W1 0_151/W2 0_110/W3 0_109/E3 0_4/N1 0_4/N2 W3 W1 x0
Xinv_customized_29 W1 0_95/W2 W3 inv_customized_29/OUT W3 W1 inv_customized
Xinv_customized_18 W1 0_157/W2 W3 inv_customized_18/OUT W3 W1 inv_customized
Xinv_customized_19 W1 0_156/W2 W3 inv_customized_19/OUT W3 W1 inv_customized
Xinv_customized_3_0 0_9/N1 W3 A2 W1 W3 W1 inv_customized_3
Xinv_customized_3_1 0_9/N2 W3 0_9/N1 W1 W3 W1 inv_customized_3
X0_90 W1 0_91/W2 0_91/W3 0_90/E3 0_9/N2 0_9/N1 W3 W1 x0
Xinv_customized_3_2 0_4/N2 W3 A1 W1 W3 W1 inv_customized_3
X0_80 W1 0_83/W2 0_81/E3 0_83/W2 0_7/N2 0_7/N1 W3 W1 x0
X0_91 W1 0_91/W2 0_91/W3 0_91/E3 0_97/N2 0_97/N1 W3 W1 x0
Xinv_customized_3_3 0_4/N1 W3 0_4/N2 W1 W3 W1 inv_customized_3
X0_70 W1 0_70/W2 W3 0_70/E3 0_79/N2 0_79/N1 W3 W1 x0
X0_81 W1 0_83/W2 0_82/E3 0_81/E3 0_4/N1 0_4/N2 W3 W1 x0
X0_92 W1 0_95/W2 0_93/W3 0_95/W2 0_7/N2 0_7/N1 W3 W1 x0
Xinv_customized_3_4 0_7/N1 W3 A0 W1 W3 W1 inv_customized_3
X0_71 W1 0_71/W2 W3 0_71/E3 0_79/N2 0_79/N1 W3 W1 x0
X0_60 W1 0_76/W2 0_60/W3 0_76/E3 0_97/N2 0_97/N1 W3 W1 x0
X0_82 W1 0_83/W2 0_83/W3 0_82/E3 0_9/N2 0_9/N1 W3 W1 x0
X0_93 W1 0_95/W2 0_93/W3 0_94/E3 0_4/N2 0_4/N1 W3 W1 x0
Xinv_customized_3_5 0_7/N2 W3 0_7/N1 W1 W3 W1 inv_customized_3
X0_72 W1 0_72/W2 W3 0_72/E3 0_79/N2 0_79/N1 W3 W1 x0
X0_61 W1 0_77/W2 0_61/W3 0_77/E3 0_97/N2 0_97/N1 W3 W1 x0
X0_50 W1 0_78/W2 0_62/W3 0_52/W3 0_9/N2 0_9/N1 W3 W1 x0
X0_83 W1 0_83/W2 0_83/W3 0_83/E3 0_97/N2 0_97/N1 W3 W1 x0
X0_94 W1 0_95/W2 0_95/W3 0_94/E3 0_9/N2 0_9/N1 W3 W1 x0
Xinv_customized_3_6 0_79/N1 W3 A4 W1 W3 W1 inv_customized_3
X0_73 W1 0_73/W2 W3 0_73/E3 0_79/N2 0_79/N1 W3 W1 x0
X0_40 W1 0_74/W2 0_40/W3 0_40/E3 0_4/N2 0_4/N1 W3 W1 x0
X0_51 W1 0_78/W2 0_78/W2 0_52/E3 0_7/N1 0_7/N2 W3 W1 x0
X0_62 W1 0_78/W2 0_62/W3 0_78/E3 0_97/N2 0_97/N1 W3 W1 x0
X0_84 W1 0_87/W2 0_87/W2 0_85/E3 0_7/N1 0_7/N2 W3 W1 x0
X0_95 W1 0_95/W2 0_95/W3 0_95/E3 0_97/N2 0_97/N1 W3 W1 x0
Xinv_customized_0 W1 0_8/W2 W3 inv_customized_0/OUT W3 W1 inv_customized
Xinv_customized_3_7 0_97/N1 W3 0_97/N2 W1 W3 W1 inv_customized_3
X0_30 W1 0_70/W2 0_70/E3 0_30/E3 0_97/N1 0_97/N2 W3 W1 x0
X0_74 W1 0_74/W2 W3 0_74/E3 0_79/N2 0_79/N1 W3 W1 x0
X0_41 W1 0_75/W2 0_43/E3 0_59/W3 0_9/N1 0_9/N2 W3 W1 x0
X0_52 W1 0_78/W2 0_52/W3 0_52/E3 0_4/N1 0_4/N2 W3 W1 x0
X0_63 W1 0_79/W2 0_63/W3 0_79/E3 0_97/N2 0_97/N1 W3 W1 x0
X0_85 W1 0_87/W2 0_86/E3 0_85/E3 0_4/N1 0_4/N2 W3 W1 x0
X0_96 W1 0_99/W2 0_99/W3 0_99/W2 0_7/N2 0_7/N1 W3 W1 x0
Xinv_customized_1 W1 0_9/W2 W3 inv_customized_1/OUT W3 W1 inv_customized
Xinv_customized_3_8 0_97/N2 W3 A3 W1 W3 W1 inv_customized_3
X0_64 W1 0_8/W2 W3 0_64/E3 0_79/N2 0_79/N1 W3 W1 x0
X0_20 W1 0_68/W2 0_20/W3 0_28/E3 0_9/N1 0_9/N2 W3 W1 x0
X0_31 W1 0_71/W2 0_71/E3 0_31/E3 0_97/N1 0_97/N2 W3 W1 x0
X0_42 W1 0_75/W2 0_43/W3 0_75/W2 0_7/N2 0_7/N1 W3 W1 x0
X0_75 W1 0_75/W2 W3 0_75/E3 0_79/N2 0_79/N1 W3 W1 x0
X0_53 W1 0_79/W2 0_54/E3 0_79/W2 0_7/N2 0_7/N1 W3 W1 x0
X0_86 W1 0_87/W2 0_87/W3 0_86/E3 0_9/N2 0_9/N1 W3 W1 x0
X0_97 W1 0_99/W2 0_98/E3 0_97/E3 0_97/N2 0_97/N1 W3 W1 x0
Xinv_customized_2 W1 0_6/W3 W3 inv_customized_2/OUT W3 W1 inv_customized
Xinv_customized_3_9 0_79/N2 W3 0_79/N1 W1 W3 W1 inv_customized_3
X0_65 W1 0_9/W2 W3 0_65/E3 0_79/N2 0_79/N1 W3 W1 x0
X0_10 W1 0_6/W3 0_26/E3 0_4/E3 0_9/N2 0_9/N1 W3 W1 x0
X0_21 W1 0_69/W2 0_21/W3 0_29/E3 0_9/N1 0_9/N2 W3 W1 x0
X0_32 W1 0_72/W2 0_34/W3 0_56/W3 0_9/N1 0_9/N2 W3 W1 x0
X0_43 W1 0_75/W2 0_43/W3 0_43/E3 0_4/N2 0_4/N1 W3 W1 x0
X0_76 W1 0_76/W2 W3 0_76/E3 0_79/N2 0_79/N1 W3 W1 x0
X0_54 W1 0_79/W2 0_55/E3 0_54/E3 0_4/N1 0_4/N2 W3 W1 x0
X0_87 W1 0_87/W2 0_87/W3 0_87/E3 0_97/N2 0_97/N1 W3 W1 x0
X0_98 W1 0_99/W2 0_99/E3 0_98/E3 0_9/N1 0_9/N2 W3 W1 x0
X0_0 W1 0_8/W2 0_8/E3 0_1/W3 0_4/N1 0_4/N2 W3 W1 x0
Xinv_customized_3 W1 0_7/W2 W3 inv_customized_3/OUT W3 W1 inv_customized
X0_66 W1 0_6/W3 W3 0_66/E3 0_79/N2 0_79/N1 W3 W1 x0
X0_11 W1 0_7/W2 0_27/E3 0_2/E3 0_9/N2 0_9/N1 W3 W1 x0
X0_22 W1 0_70/W2 0_22/W3 0_30/E3 0_9/N1 0_9/N2 W3 W1 x0
X0_33 W1 0_72/W2 0_34/E3 0_72/W2 0_7/N2 0_7/N1 W3 W1 x0
X0_44 W1 0_76/W2 0_60/W3 0_46/E3 0_9/N2 0_9/N1 W3 W1 x0
X0_55 W1 0_79/W2 0_63/W3 0_55/E3 0_9/N2 0_9/N1 W3 W1 x0
X0_1 W1 0_8/W2 0_1/W3 0_8/W2 0_7/N2 0_7/N1 W3 W1 x0
X0_77 W1 0_77/W2 W3 0_77/E3 0_79/N2 0_79/N1 W3 W1 x0
X0_88 W1 0_91/W2 0_91/W2 0_89/W3 0_7/N1 0_7/N2 W3 W1 x0
X0_99 W1 0_99/W2 0_99/W3 0_99/E3 0_4/N2 0_4/N1 W3 W1 x0
Xinv_customized_4 W1 0_68/W2 W3 inv_customized_4/OUT W3 W1 inv_customized
X0_67 W1 0_7/W2 W3 0_67/E3 0_79/N2 0_79/N1 W3 W1 x0
X0_12 W1 0_68/W2 0_13/W3 0_20/W3 0_4/N2 0_4/N1 W3 W1 x0
X0_23 W1 0_71/W2 0_23/W3 0_31/E3 0_9/N1 0_9/N2 W3 W1 x0
X0_34 W1 0_72/W2 0_34/W3 0_34/E3 0_4/N1 0_4/N2 W3 W1 x0
X0_56 W1 0_72/W2 0_56/W3 0_72/E3 0_97/N2 0_97/N1 W3 W1 x0
X0_45 W1 0_76/W2 0_46/W3 0_76/W2 0_7/N2 0_7/N1 W3 W1 x0
X0_78 W1 0_78/W2 W3 0_78/E3 0_79/N2 0_79/N1 W3 W1 x0
X0_89 W1 0_91/W2 0_89/W3 0_90/E3 0_4/N2 0_4/N1 W3 W1 x0
X0_2 W1 0_7/W2 0_7/W3 0_2/E3 0_4/N2 0_4/N1 W3 W1 x0
Xinv_customized_5 W1 0_69/W2 W3 inv_customized_5/OUT W3 W1 inv_customized
X0_24 W1 0_8/W2 0_64/E3 0_8/W3 0_97/N1 0_97/N2 W3 W1 x0
X0_3 W1 0_9/W2 0_9/E3 0_5/E3 0_4/N1 0_4/N2 W3 W1 x0
X0_13 W1 0_68/W2 0_13/W3 0_68/W2 0_7/N2 0_7/N1 W3 W1 x0
X0_68 W1 0_68/W2 W3 0_68/E3 0_79/N2 0_79/N1 W3 W1 x0
X0_35 W1 0_73/W2 0_37/W3 0_57/W3 0_9/N1 0_9/N2 W3 W1 x0
X0_57 W1 0_73/W2 0_57/W3 0_73/E3 0_97/N2 0_97/N1 W3 W1 x0
X0_46 W1 0_76/W2 0_46/W3 0_46/E3 0_4/N2 0_4/N1 W3 W1 x0
X0_79 W1 0_79/W2 W3 0_79/E3 0_79/N2 0_79/N1 W3 W1 x0
Xinv_customized_6 W1 0_70/W2 W3 inv_customized_6/OUT W3 W1 inv_customized
X0_25 W1 0_9/W2 0_65/E3 0_9/W3 0_97/N1 0_97/N2 W3 W1 x0
X0_14 W1 0_69/W2 0_69/W2 0_15/W3 0_7/N1 0_7/N2 W3 W1 x0
X0_69 W1 0_69/W2 W3 0_69/E3 0_79/N2 0_79/N1 W3 W1 x0
X0_36 W1 0_73/W2 0_73/W2 0_37/E3 0_7/N1 0_7/N2 W3 W1 x0
X0_58 W1 0_74/W2 0_58/W3 0_74/E3 0_97/N2 0_97/N1 W3 W1 x0
X0_47 W1 0_77/W2 0_61/W3 0_49/E3 0_9/N2 0_9/N1 W3 W1 x0
X0_4 W1 0_6/W3 0_6/E3 0_4/E3 0_4/N2 0_4/N1 W3 W1 x0
Xinv_customized_7 W1 0_71/W2 W3 inv_customized_7/OUT W3 W1 inv_customized
X0_5 W1 0_9/W2 0_9/W2 0_5/E3 0_7/N1 0_7/N2 W3 W1 x0
X0_26 W1 0_6/W3 0_66/E3 0_26/E3 0_97/N1 0_97/N2 W3 W1 x0
X0_15 W1 0_69/W2 0_15/W3 0_21/W3 0_4/N2 0_4/N1 W3 W1 x0
X0_37 W1 0_73/W2 0_37/W3 0_37/E3 0_4/N1 0_4/N2 W3 W1 x0
X0_59 W1 0_75/W2 0_59/W3 0_75/E3 0_97/N2 0_97/N1 W3 W1 x0
X0_48 W1 0_77/W2 0_77/W2 0_49/W3 0_7/N1 0_7/N2 W3 W1 x0
X0_150 W1 0_150/W2 0_150/W3 W3 0_79/N1 0_79/N2 W3 W1 x0
Xinv_customized_8 W1 0_78/W2 W3 inv_customized_8/OUT W3 W1 inv_customized
X0_27 W1 0_7/W2 0_67/E3 0_27/E3 0_97/N1 0_97/N2 W3 W1 x0
X0_16 W1 0_70/W2 0_22/W3 0_17/E3 0_4/N1 0_4/N2 W3 W1 x0
X0_38 W1 0_74/W2 0_40/E3 0_58/W3 0_9/N1 0_9/N2 W3 W1 x0
X0_49 W1 0_77/W2 0_49/W3 0_49/E3 0_4/N2 0_4/N1 W3 W1 x0
X0_6 W1 0_6/W3 0_6/W3 0_6/E3 0_7/N1 0_7/N2 W3 W1 x0
X0_140 W1 0_159/W2 0_141/E3 0_159/W2 0_7/N2 0_7/N1 W3 W1 x0
X0_151 W1 0_151/W2 0_151/W3 W3 0_79/N1 0_79/N2 W3 W1 x0
Xinv_customized_9 W1 0_77/W2 W3 inv_customized_9/OUT W3 W1 inv_customized
X0_7 W1 0_7/W2 0_7/W3 0_7/W2 0_7/N2 0_7/N1 W3 W1 x0
X0_28 W1 0_68/W2 0_68/E3 0_28/E3 0_97/N1 0_97/N2 W3 W1 x0
X0_17 W1 0_70/W2 0_70/W2 0_17/E3 0_7/N1 0_7/N2 W3 W1 x0
X0_39 W1 0_74/W2 0_74/W2 0_40/W3 0_7/N1 0_7/N2 W3 W1 x0
X0_141 W1 0_159/W2 0_142/E3 0_141/E3 0_4/N1 0_4/N2 W3 W1 x0
X0_130 W1 0_156/W2 0_156/W3 0_130/E3 0_97/N1 0_97/N2 W3 W1 x0
X0_152 W1 0_152/W2 0_152/W3 W3 0_79/N1 0_79/N2 W3 W1 x0
X0_29 W1 0_69/W2 0_69/E3 0_29/E3 0_97/N1 0_97/N2 W3 W1 x0
X0_18 W1 0_71/W2 0_23/W3 0_19/W3 0_4/N1 0_4/N2 W3 W1 x0
X0_8 W1 0_8/W2 0_8/W3 0_8/E3 0_9/N2 0_9/N1 W3 W1 x0
X0_142 W1 0_159/W2 0_143/E3 0_142/E3 0_9/N2 0_9/N1 W3 W1 x0
X0_131 W1 0_156/W2 0_131/W3 0_131/E3 0_4/N2 0_4/N1 W3 W1 x0
X0_120 W1 0_154/W2 0_154/W2 0_123/W3 0_7/N1 0_7/N2 W3 W1 x0
X0_153 W1 0_153/W2 0_153/W3 W3 0_79/N1 0_79/N2 W3 W1 x0
X0_19 W1 0_71/W2 0_19/W3 0_71/W2 0_7/N2 0_7/N1 W3 W1 x0
X0_9 W1 0_9/W2 0_9/W3 0_9/E3 0_9/N2 0_9/N1 W3 W1 x0
X0_143 W1 0_159/W2 0_159/W3 0_143/E3 0_97/N1 0_97/N2 W3 W1 x0
X0_132 W1 0_157/W2 0_157/W2 0_135/W3 0_7/N1 0_7/N2 W3 W1 x0
X0_121 W1 0_154/W2 0_154/W3 0_122/E3 0_97/N1 0_97/N2 W3 W1 x0
X0_154 W1 0_154/W2 0_154/W3 W3 0_79/N1 0_79/N2 W3 W1 x0
X0_110 W1 0_151/W2 0_110/W3 0_111/W3 0_9/N1 0_9/N2 W3 W1 x0
Xinv_customized_30 W1 0_87/W2 W3 inv_customized_30/OUT W3 W1 inv_customized
X0_144 W1 0_83/W2 0_83/E3 W3 0_79/N1 0_79/N2 W3 W1 x0
X0_133 W1 0_157/W2 0_157/W3 0_134/W3 0_97/N1 0_97/N2 W3 W1 x0
X0_155 W1 0_155/W2 0_155/W3 W3 0_79/N1 0_79/N2 W3 W1 x0
X0_122 W1 0_154/W2 0_123/E3 0_122/E3 0_9/N1 0_9/N2 W3 W1 x0
X0_111 W1 0_151/W2 0_111/W3 0_151/W3 0_97/N2 0_97/N1 W3 W1 x0
X0_100 W1 0_149/W2 0_149/W2 0_101/W3 0_7/N1 0_7/N2 W3 W1 x0
Xinv_customized_31 W1 0_83/W2 W3 inv_customized_31/OUT W3 W1 inv_customized
Xinv_customized_20 W1 0_155/W2 W3 inv_customized_20/OUT W3 W1 inv_customized
X0_145 W1 0_87/W2 0_87/E3 W3 0_79/N1 0_79/N2 W3 W1 x0
X0_134 W1 0_157/W2 0_134/W3 0_135/E3 0_9/N2 0_9/N1 W3 W1 x0
X0_156 W1 0_156/W2 0_156/W3 W3 0_79/N1 0_79/N2 W3 W1 x0
X0_123 W1 0_154/W2 0_123/W3 0_123/E3 0_4/N2 0_4/N1 W3 W1 x0
X0_112 W1 0_152/W2 0_115/E3 0_152/W2 0_7/N2 0_7/N1 W3 W1 x0
X0_101 W1 0_149/W2 0_101/W3 0_102/W3 0_4/N2 0_4/N1 W3 W1 x0
Xinv_customized_10 W1 0_76/W2 W3 inv_customized_10/OUT W3 W1 inv_customized
Xinv_customized_21 W1 0_154/W2 W3 inv_customized_21/OUT W3 W1 inv_customized
X0_146 W1 0_91/W2 0_91/E3 W3 0_79/N1 0_79/N2 W3 W1 x0
X0_157 W1 0_157/W2 0_157/W3 W3 0_79/N1 0_79/N2 W3 W1 x0
X0_135 W1 0_157/W2 0_135/W3 0_135/E3 0_4/N2 0_4/N1 W3 W1 x0
X0_124 W1 0_155/W2 0_125/W3 0_155/W2 0_7/N2 0_7/N1 W3 W1 x0
X0_113 W1 0_152/W2 0_152/W3 0_114/E3 0_97/N1 0_97/N2 W3 W1 x0
X0_102 W1 0_149/W2 0_102/W3 0_103/W3 0_9/N1 0_9/N2 W3 W1 x0
Xinv_customized_11 W1 0_75/W2 W3 inv_customized_11/OUT W3 W1 inv_customized
Xinv_customized_22 W1 0_153/W2 W3 inv_customized_22/OUT W3 W1 inv_customized
X0_147 W1 0_95/W2 0_95/E3 W3 0_79/N1 0_79/N2 W3 W1 x0
X0_158 W1 0_158/W2 0_158/W3 W3 0_79/N1 0_79/N2 W3 W1 x0
X0_136 W1 0_158/W2 0_158/W2 0_137/E3 0_7/N1 0_7/N2 W3 W1 x0
X0_125 W1 0_155/W2 0_125/W3 0_126/W3 0_4/N2 0_4/N1 W3 W1 x0
X0_114 W1 0_152/W2 0_115/W3 0_114/E3 0_9/N1 0_9/N2 W3 W1 x0
X0_103 W1 0_149/W2 0_103/W3 0_149/W3 0_97/N2 0_97/N1 W3 W1 x0
Xinv_customized_12 W1 0_74/W2 W3 inv_customized_12/OUT W3 W1 inv_customized
Xinv_customized_23 W1 0_152/W2 W3 inv_customized_23/OUT W3 W1 inv_customized
X0_148 W1 0_99/W2 0_97/E3 W3 0_79/N1 0_79/N2 W3 W1 x0
X0_159 W1 0_159/W2 0_159/W3 W3 0_79/N1 0_79/N2 W3 W1 x0
X0_137 W1 0_158/W2 0_138/E3 0_137/E3 0_4/N1 0_4/N2 W3 W1 x0
X0_126 W1 0_155/W2 0_126/W3 0_127/E3 0_9/N1 0_9/N2 W3 W1 x0
X0_115 W1 0_152/W2 0_115/W3 0_115/E3 0_4/N1 0_4/N2 W3 W1 x0
X0_104 W1 0_150/W2 0_150/W2 0_105/E3 0_7/N1 0_7/N2 W3 W1 x0
Xinv_customized_13 W1 0_73/W2 W3 inv_customized_13/OUT W3 W1 inv_customized
Xinv_customized_24 W1 0_150/W2 W3 inv_customized_24/OUT W3 W1 inv_customized
C0 0_4/N2 W1 2.03fF
C1 W1 W3 167.25fF
C2 0_159/W2 W3 2.98fF
C3 0_99/W2 W3 3.02fF
C4 0_158/W2 W3 2.87fF
C5 0_95/W2 W3 2.93fF
C6 0_157/W2 W3 2.83fF
C7 0_91/W2 W3 2.88fF
C8 0_156/W2 W3 3.01fF
C9 0_87/W2 W3 2.83fF
C10 0_155/W2 W3 2.93fF
C11 0_83/W2 W3 3.03fF
C12 0_154/W2 W3 2.88fF
C13 0_153/W2 W3 2.83fF
C14 0_152/W2 W3 3.02fF
C15 0_151/W2 W3 2.93fF
C16 0_150/W2 W3 2.88fF
C17 0_69/W2 W3 2.83fF
C18 0_79/W2 W3 2.93fF
C19 0_68/W2 W3 2.98fF
C20 0_78/W2 W3 2.87fF
C21 0_7/W2 W3 2.93fF
C22 0_77/W2 W3 2.83fF
C23 0_6/W3 W3 2.88fF
C24 0_76/W2 W3 3.01fF
C25 0_9/W2 W3 2.83fF
C26 0_79/N2 W3 24.71fF
C27 0_79/N1 W3 24.32fF
C28 0_75/W2 W3 2.93fF
C29 0_8/W2 W3 2.99fF
C30 0_97/N2 W3 24.69fF
C31 0_74/W2 W3 2.87fF
C32 0_97/N1 W3 24.73fF
C33 0_73/W2 W3 2.83fF
C34 0_72/W2 W3 2.98fF
C35 0_7/N2 W3 21.79fF
C36 0_7/N1 W3 21.17fF
C37 0_71/W2 W3 2.93fF
C38 0_70/W2 W3 2.88fF
C39 0_4/N1 W3 21.88fF
C40 0_4/N2 W3 22.07fF
C41 0_9/N2 W3 15.45fF
C42 0_9/N1 W3 23.87fF
C43 0_149/W2 W3 2.83fF
.ends

