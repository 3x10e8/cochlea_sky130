magic
tech sky130A
timestamp 1639199554
<< nwell >>
rect 106 301 262 519
<< nmos >>
rect 175 142 193 242
<< pmos >>
rect 175 360 193 460
<< ndiff >>
rect 125 229 175 242
rect 125 211 142 229
rect 159 211 175 229
rect 125 173 175 211
rect 125 155 142 173
rect 159 155 175 173
rect 125 142 175 155
rect 193 229 243 242
rect 193 211 209 229
rect 226 211 243 229
rect 193 173 243 211
rect 193 155 209 173
rect 226 155 243 173
rect 193 142 243 155
<< pdiff >>
rect 125 447 175 460
rect 125 429 142 447
rect 159 429 175 447
rect 125 391 175 429
rect 125 373 142 391
rect 159 373 175 391
rect 125 360 175 373
rect 193 447 243 460
rect 193 429 209 447
rect 226 429 243 447
rect 193 391 243 429
rect 193 373 209 391
rect 226 373 243 391
rect 193 360 243 373
<< ndiffc >>
rect 142 211 159 229
rect 142 155 159 173
rect 209 211 226 229
rect 209 155 226 173
<< pdiffc >>
rect 142 429 159 447
rect 142 373 159 391
rect 209 429 226 447
rect 209 373 226 391
<< poly >>
rect 167 502 201 510
rect 167 484 175 502
rect 193 484 201 502
rect 167 474 201 484
rect 175 460 193 474
rect 175 346 193 360
rect 167 336 201 346
rect 167 318 175 336
rect 193 318 201 336
rect 167 282 201 318
rect 167 264 175 282
rect 193 264 201 282
rect 167 256 201 264
rect 175 242 193 256
rect 175 128 193 142
rect 167 120 201 128
rect 167 102 175 120
rect 193 102 201 120
rect 167 94 201 102
<< polycont >>
rect 175 484 193 502
rect 175 318 193 336
rect 175 264 193 282
rect 175 102 193 120
<< locali >>
rect 167 509 201 510
rect 167 482 169 509
rect 199 482 201 509
rect 167 474 201 482
rect 132 447 168 456
rect 132 429 142 447
rect 159 429 168 447
rect 132 420 168 429
rect 200 450 236 456
rect 231 423 236 450
rect 200 420 236 423
rect 132 395 168 400
rect 163 368 168 395
rect 132 364 168 368
rect 200 391 236 400
rect 200 373 209 391
rect 226 373 236 391
rect 200 364 236 373
rect 167 336 201 346
rect 167 318 175 336
rect 193 318 201 336
rect 167 317 201 318
rect 167 290 169 317
rect 199 290 201 317
rect 167 282 201 290
rect 167 264 175 282
rect 193 264 201 282
rect 167 256 201 264
rect 132 229 168 238
rect 132 211 142 229
rect 159 211 168 229
rect 132 202 168 211
rect 200 229 236 238
rect 200 211 209 229
rect 226 211 236 229
rect 200 202 236 211
rect 132 178 168 182
rect 163 151 168 178
rect 132 146 168 151
rect 200 178 236 182
rect 200 151 204 178
rect 235 151 236 178
rect 200 146 236 151
rect 167 122 201 128
rect 167 95 169 122
rect 199 95 201 122
rect 167 94 201 95
<< viali >>
rect 169 502 199 509
rect 169 484 175 502
rect 175 484 193 502
rect 193 484 199 502
rect 169 482 199 484
rect 200 447 231 450
rect 200 429 209 447
rect 209 429 226 447
rect 226 429 231 447
rect 200 423 231 429
rect 132 391 163 395
rect 132 373 142 391
rect 142 373 159 391
rect 159 373 163 391
rect 132 368 163 373
rect 169 290 199 317
rect 132 173 163 178
rect 132 155 142 173
rect 142 155 159 173
rect 159 155 163 173
rect 132 151 163 155
rect 204 173 235 178
rect 204 155 209 173
rect 209 155 226 173
rect 226 155 235 173
rect 204 151 235 155
rect 169 120 199 122
rect 169 102 175 120
rect 175 102 193 120
rect 193 102 199 120
rect 169 95 199 102
<< metal1 >>
rect 162 509 205 514
rect 162 482 169 509
rect 199 482 205 509
rect 162 475 205 482
rect 195 454 252 459
rect -88 450 334 454
rect -88 426 200 450
rect 195 423 200 426
rect 231 426 334 450
rect 231 423 252 426
rect 195 416 252 423
rect 111 395 168 402
rect 111 387 132 395
rect -89 368 132 387
rect 163 387 168 395
rect 163 368 335 387
rect -89 359 335 368
rect 162 317 205 322
rect 162 290 169 317
rect 199 290 205 317
rect 162 283 205 290
rect 112 178 169 185
rect 112 170 132 178
rect -88 151 132 170
rect 163 151 169 178
rect -88 142 169 151
rect 199 178 256 184
rect 199 151 204 178
rect 235 171 256 178
rect 235 151 335 171
rect 199 142 335 151
rect 199 141 256 142
rect 162 122 205 127
rect 162 95 169 122
rect 199 95 205 122
rect 162 88 205 95
<< via1 >>
rect 169 482 199 509
rect 169 290 199 317
rect 169 95 199 122
<< metal2 >>
rect 40 47 84 560
rect 162 509 205 561
rect 162 482 169 509
rect 199 482 205 509
rect 162 475 205 482
rect 162 317 205 322
rect 162 290 169 317
rect 199 290 205 317
rect 162 283 205 290
rect 162 122 205 127
rect 162 95 169 122
rect 199 95 205 122
rect 162 48 205 95
<< labels >>
rlabel metal2 186 560 186 560 1 N1
port 9 n
rlabel metal2 61 559 61 559 1 N2
port 10 n
rlabel metal1 333 440 333 440 3 W1
port 8 e
rlabel metal1 334 371 334 371 3 W2
port 7 e
rlabel metal1 334 156 334 156 3 W3
port 6 e
rlabel metal1 -87 440 -87 440 7 E1
port 1 w
rlabel metal1 -88 373 -88 373 7 E2
port 2 w
rlabel metal1 -87 157 -87 157 7 E3
port 3 w
rlabel metal2 63 48 63 48 5 S2
port 4 s
rlabel metal2 185 49 185 49 5 S1
port 5 s
<< end >>
