* SPICE3 file created from /home/sky/Desktop/BENG207_Project/cochlea_sky130/mag/HW4_layout/2x4/2x4_circuit.ext - technology: sky130A

.subckt x1 W1 W2 E3 S2 S1 W3 SUB
X0 W1 S1 W2 w_106_301# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X1 W3 S1 E3 SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
.ends

.subckt inv_customized GND IN VDD SUB OUT
X0 OUT IN VDD w_n16_301# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X1 OUT IN GND SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
.ends

.subckt x0_unit W3 S1 S2 E3 W2 W1 SUB
X0 W2 S1 W1 w_n16_301# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X1 E3 S1 W3 SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
.ends

.subckt x/home/sky/Desktop/BENG207_Project/cochlea_sky130/mag/HW4_layout/2x4/2x4_circuit
+ Gate
X1_0 W1 1_0/W3 1_0/E3 1_1/S2 1_1/S1 1_0/W3 SUB x1
X1_1 W1 1_2/W2 1_2/W3 1_1/S2 1_1/S1 1_2/W2 SUB x1
X1_2 W1 1_2/W2 W3 Gate S2 1_2/W3 SUB x1
X1_3 W1 1_3/W2 W3 Gate S2 1_3/W3 SUB x1
Xinv_customized_0 W3 W2 W1 SUB sel0 inv_customized
Xinv_customized_1 W3 1_0/W3 W1 SUB sel1 inv_customized
X0_unit_0 E3 1_1/S2 1_1/S1 W2 W2 W1 SUB x0_unit
Xinv_customized_2 W3 1_2/W2 W1 SUB sel2 inv_customized
X0_unit_1 W3 Gate S2 1_0/E3 1_0/W3 W1 SUB x0_unit
Xinv_customized_3 W3 1_3/W2 W1 SUB sel3 inv_customized
Xinv_customized_4 W3 1_1/S2 W1 SUB 1_1/S1 inv_customized
X0_unit_2 1_3/W3 1_1/S2 1_1/S1 1_3/W2 1_3/W2 W1 SUB x0_unit
Xinv_customized_5 W3 Gate W1 SUB S2 inv_customized
Xinv_customized_6 W3 A1 W1 SUB Gate inv_customized
Xinv_customized_7 W3 A0 W1 SUB 1_1/S2 inv_customized
X0 W2 Gate W1 w_n16_301# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X1 E3 Gate W3 SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
C0 W3 Gate 2.03fF
C1 W3 SUB -4.59fF
C2 W1 SUB -6.10fF
C3 1_1/S1 SUB 2.34fF
C4 1_1/S2 SUB 4.86fF
C5 S2 SUB 2.25fF
.ends

