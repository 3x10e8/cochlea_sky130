magic
tech sky130A
timestamp 1639220931
<< nwell >>
rect 2067 283 4452 439
rect 2067 -229 4452 -73
rect 2067 -758 4452 -602
rect 2067 -1280 4452 -1124
rect 2065 -1806 4450 -1650
rect 2067 -2330 4452 -2174
rect 2067 -2854 4452 -2698
rect 2063 -3372 4448 -3216
rect 2065 -3901 4450 -3745
rect 2067 -4419 4452 -4263
rect 2065 -4947 4450 -4791
rect 2067 -5469 4452 -5313
rect 2067 -5985 4452 -5829
rect 2067 -6510 4452 -6354
rect 2067 -7034 4452 -6878
rect 2067 -7558 4452 -7402
rect 2189 -8076 4449 -7923
rect 2189 -8603 4449 -8450
rect 2189 -9122 4449 -8969
rect 2187 -9647 4447 -9494
rect 2189 -10164 4449 -10011
rect 2189 -10687 4449 -10534
rect 2189 -11214 4449 -11061
rect 2189 -11733 4449 -11580
rect 2189 -12260 4449 -12107
rect 2189 -12787 4449 -12634
rect 2189 -13307 4449 -13154
rect 2189 -13828 4449 -13675
rect 2189 -14348 4449 -14195
rect 2189 -14872 4449 -14719
rect 2189 -15395 4449 -15242
rect 2185 -15908 4445 -15755
rect 2074 -16919 2187 -16520
rect 2507 -16925 2620 -16526
rect 2929 -16923 3042 -16524
rect 3355 -16925 3468 -16526
rect 3777 -16927 3890 -16528
<< metal1 >>
rect 1534 360 1826 508
rect 1534 305 2029 360
rect 1534 -163 1826 305
rect 1887 78 1979 83
rect 1887 0 1892 78
rect 1970 72 1979 78
rect 1970 11 2037 72
rect 1970 0 1979 11
rect 1887 -9 1979 0
rect 1534 -218 2029 -163
rect 1534 -686 1826 -218
rect 1887 -445 1979 -440
rect 1887 -523 1892 -445
rect 1970 -451 1979 -445
rect 1970 -512 2037 -451
rect 1970 -523 1979 -512
rect 1887 -532 1979 -523
rect 1534 -741 2029 -686
rect 1534 -1209 1826 -741
rect 1887 -968 1979 -963
rect 1887 -1046 1892 -968
rect 1970 -974 1979 -968
rect 1970 -1035 2037 -974
rect 1970 -1046 1979 -1035
rect 1887 -1055 1979 -1046
rect 1534 -1264 2029 -1209
rect 1534 -1732 1826 -1264
rect 1887 -1491 1979 -1486
rect 1887 -1569 1892 -1491
rect 1970 -1497 1979 -1491
rect 1970 -1558 2037 -1497
rect 1970 -1569 1979 -1558
rect 1887 -1578 1979 -1569
rect 1534 -1787 2029 -1732
rect 1534 -2255 1826 -1787
rect 1887 -2014 1979 -2009
rect 1887 -2092 1892 -2014
rect 1970 -2020 1979 -2014
rect 1970 -2081 2037 -2020
rect 1970 -2092 1979 -2081
rect 1887 -2101 1979 -2092
rect 1534 -2310 2029 -2255
rect 1534 -2778 1826 -2310
rect 1887 -2537 1979 -2532
rect 1887 -2615 1892 -2537
rect 1970 -2543 1979 -2537
rect 1970 -2604 2037 -2543
rect 1970 -2615 1979 -2604
rect 1887 -2624 1979 -2615
rect 1534 -2833 2029 -2778
rect 1534 -3301 1826 -2833
rect 1887 -3060 1979 -3055
rect 1887 -3138 1892 -3060
rect 1970 -3066 1979 -3060
rect 1970 -3127 2037 -3066
rect 1970 -3138 1979 -3127
rect 1887 -3147 1979 -3138
rect 1534 -3356 2029 -3301
rect 1534 -3824 1826 -3356
rect 1887 -3583 1979 -3578
rect 1887 -3661 1892 -3583
rect 1970 -3589 1979 -3583
rect 1970 -3650 2037 -3589
rect 1970 -3661 1979 -3650
rect 1887 -3670 1979 -3661
rect 1534 -3879 2029 -3824
rect 1534 -4347 1826 -3879
rect 1887 -4106 1979 -4101
rect 1887 -4184 1892 -4106
rect 1970 -4112 1979 -4106
rect 1970 -4173 2037 -4112
rect 1970 -4184 1979 -4173
rect 1887 -4193 1979 -4184
rect 1534 -4402 2029 -4347
rect 1534 -4870 1826 -4402
rect 1887 -4629 1979 -4624
rect 1887 -4707 1892 -4629
rect 1970 -4635 1979 -4629
rect 1970 -4696 2037 -4635
rect 1970 -4707 1979 -4696
rect 1887 -4716 1979 -4707
rect 1534 -4925 2029 -4870
rect 1534 -5393 1826 -4925
rect 1887 -5152 1979 -5147
rect 1887 -5230 1892 -5152
rect 1970 -5158 1979 -5152
rect 1970 -5219 2037 -5158
rect 1970 -5230 1979 -5219
rect 1887 -5239 1979 -5230
rect 1534 -5448 2029 -5393
rect 1534 -5916 1826 -5448
rect 1887 -5675 1979 -5670
rect 1887 -5753 1892 -5675
rect 1970 -5681 1979 -5675
rect 1970 -5742 2037 -5681
rect 1970 -5753 1979 -5742
rect 1887 -5762 1979 -5753
rect 1534 -5971 2029 -5916
rect 1534 -6439 1826 -5971
rect 1887 -6198 1979 -6193
rect 1887 -6276 1892 -6198
rect 1970 -6204 1979 -6198
rect 1970 -6265 2037 -6204
rect 1970 -6276 1979 -6265
rect 1887 -6285 1979 -6276
rect 1534 -6494 2029 -6439
rect 1534 -6962 1826 -6494
rect 1887 -6721 1979 -6716
rect 1887 -6799 1892 -6721
rect 1970 -6727 1979 -6721
rect 1970 -6788 2037 -6727
rect 1970 -6799 1979 -6788
rect 1887 -6808 1979 -6799
rect 1534 -7017 2029 -6962
rect 1534 -7485 1826 -7017
rect 1887 -7244 1979 -7239
rect 1887 -7322 1892 -7244
rect 1970 -7250 1979 -7244
rect 1970 -7311 2037 -7250
rect 1970 -7322 1979 -7311
rect 1887 -7331 1979 -7322
rect 1534 -7540 2029 -7485
rect 1534 -8008 1826 -7540
rect 1887 -7767 1979 -7762
rect 1887 -7845 1892 -7767
rect 1970 -7773 1979 -7767
rect 1970 -7834 2037 -7773
rect 1970 -7845 1979 -7834
rect 1887 -7854 1979 -7845
rect 1534 -8063 2029 -8008
rect 1534 -8531 1826 -8063
rect 1887 -8290 1979 -8285
rect 1887 -8368 1892 -8290
rect 1970 -8296 1979 -8290
rect 1970 -8357 2037 -8296
rect 1970 -8368 1979 -8357
rect 1887 -8377 1979 -8368
rect 1534 -8586 2029 -8531
rect 1534 -9054 1826 -8586
rect 1887 -8813 1979 -8808
rect 1887 -8891 1892 -8813
rect 1970 -8819 1979 -8813
rect 1970 -8880 2037 -8819
rect 1970 -8891 1979 -8880
rect 1887 -8900 1979 -8891
rect 1534 -9109 2029 -9054
rect 1534 -9577 1826 -9109
rect 1887 -9336 1979 -9331
rect 1887 -9414 1892 -9336
rect 1970 -9342 1979 -9336
rect 1970 -9403 2037 -9342
rect 1970 -9414 1979 -9403
rect 1887 -9423 1979 -9414
rect 1534 -9632 2029 -9577
rect 1534 -10100 1826 -9632
rect 1887 -9859 1979 -9854
rect 1887 -9937 1892 -9859
rect 1970 -9865 1979 -9859
rect 1970 -9926 2037 -9865
rect 1970 -9937 1979 -9926
rect 1887 -9946 1979 -9937
rect 1534 -10155 2029 -10100
rect 1534 -10623 1826 -10155
rect 1887 -10382 1979 -10377
rect 1887 -10460 1892 -10382
rect 1970 -10388 1979 -10382
rect 1970 -10449 2037 -10388
rect 1970 -10460 1979 -10449
rect 1887 -10469 1979 -10460
rect 1534 -10678 2029 -10623
rect 1534 -11146 1826 -10678
rect 1887 -10905 1979 -10900
rect 1887 -10983 1892 -10905
rect 1970 -10911 1979 -10905
rect 1970 -10972 2037 -10911
rect 1970 -10983 1979 -10972
rect 1887 -10992 1979 -10983
rect 1534 -11201 2029 -11146
rect 1534 -11669 1826 -11201
rect 1887 -11428 1979 -11423
rect 1887 -11506 1892 -11428
rect 1970 -11434 1979 -11428
rect 1970 -11495 2037 -11434
rect 1970 -11506 1979 -11495
rect 1887 -11515 1979 -11506
rect 1534 -11724 2029 -11669
rect 1534 -12192 1826 -11724
rect 1887 -11951 1979 -11946
rect 1887 -12029 1892 -11951
rect 1970 -11957 1979 -11951
rect 1970 -12018 2037 -11957
rect 1970 -12029 1979 -12018
rect 1887 -12038 1979 -12029
rect 1534 -12247 2029 -12192
rect 1534 -12715 1826 -12247
rect 1887 -12474 1979 -12469
rect 1887 -12552 1892 -12474
rect 1970 -12480 1979 -12474
rect 1970 -12541 2037 -12480
rect 1970 -12552 1979 -12541
rect 1887 -12561 1979 -12552
rect 1534 -12770 2029 -12715
rect 1534 -13238 1826 -12770
rect 1887 -12997 1979 -12992
rect 1887 -13075 1892 -12997
rect 1970 -13003 1979 -12997
rect 1970 -13064 2037 -13003
rect 1970 -13075 1979 -13064
rect 1887 -13084 1979 -13075
rect 1534 -13293 2029 -13238
rect 1534 -13761 1826 -13293
rect 1887 -13520 1979 -13515
rect 1887 -13598 1892 -13520
rect 1970 -13526 1979 -13520
rect 1970 -13587 2037 -13526
rect 1970 -13598 1979 -13587
rect 1887 -13607 1979 -13598
rect 1534 -13816 2029 -13761
rect 1534 -14284 1826 -13816
rect 1887 -14043 1979 -14038
rect 1887 -14121 1892 -14043
rect 1970 -14049 1979 -14043
rect 1970 -14110 2037 -14049
rect 1970 -14121 1979 -14110
rect 1887 -14130 1979 -14121
rect 1534 -14339 2029 -14284
rect 1534 -14807 1826 -14339
rect 1887 -14566 1979 -14561
rect 1887 -14644 1892 -14566
rect 1970 -14572 1979 -14566
rect 1970 -14633 2037 -14572
rect 1970 -14644 1979 -14633
rect 1887 -14653 1979 -14644
rect 1534 -14862 2029 -14807
rect 1534 -15330 1826 -14862
rect 1887 -15089 1979 -15084
rect 1887 -15167 1892 -15089
rect 1970 -15095 1979 -15089
rect 1970 -15156 2037 -15095
rect 1970 -15167 1979 -15156
rect 1887 -15176 1979 -15167
rect 1534 -15385 2029 -15330
rect 1534 -15853 1826 -15385
rect 1887 -15612 1979 -15607
rect 1887 -15690 1892 -15612
rect 1970 -15618 1979 -15612
rect 1970 -15679 2037 -15618
rect 1970 -15690 1979 -15679
rect 1887 -15699 1979 -15690
rect 1534 -15908 2029 -15853
rect 1534 -16629 1826 -15908
rect 1947 -16125 2039 -16116
rect 1947 -16208 1956 -16125
rect 2029 -16208 2039 -16125
rect 1947 -16217 2039 -16208
rect 2653 -16301 2729 -16300
rect 2231 -16308 2304 -16306
rect 2231 -16356 2236 -16308
rect 2301 -16356 2304 -16308
rect 2231 -16363 2304 -16356
rect 2653 -16350 2658 -16301
rect 2725 -16350 2729 -16301
rect 2653 -16358 2729 -16350
rect 3080 -16304 3153 -16301
rect 3929 -16304 4002 -16301
rect 3080 -16352 3083 -16304
rect 3148 -16352 3153 -16304
rect 3080 -16358 3153 -16352
rect 3506 -16308 3579 -16304
rect 3506 -16356 3511 -16308
rect 3576 -16356 3579 -16308
rect 3506 -16361 3579 -16356
rect 3929 -16352 3932 -16304
rect 3997 -16352 4002 -16304
rect 3929 -16358 4002 -16352
rect 2098 -16629 2123 -16540
rect 2640 -16549 2716 -16545
rect 2523 -16629 2550 -16555
rect 2640 -16598 2645 -16549
rect 2712 -16598 2716 -16549
rect 2640 -16603 2716 -16598
rect 2949 -16629 2974 -16549
rect 3375 -16629 3400 -16538
rect 3803 -16629 3825 -16498
rect 1534 -16679 4201 -16629
rect 1534 -17023 1826 -16679
rect 2523 -16696 2550 -16679
rect 2949 -16680 2974 -16679
rect 3078 -16702 3151 -16700
rect 2229 -16707 2302 -16702
rect 2229 -16755 2233 -16707
rect 2298 -16755 2302 -16707
rect 2229 -16759 2302 -16755
rect 2653 -16706 2729 -16702
rect 2653 -16755 2656 -16706
rect 2723 -16755 2729 -16706
rect 2653 -16760 2729 -16755
rect 3078 -16750 3083 -16702
rect 3148 -16750 3151 -16702
rect 3078 -16757 3151 -16750
rect 3502 -16704 3575 -16700
rect 3502 -16752 3506 -16704
rect 3571 -16752 3575 -16704
rect 3502 -16757 3575 -16752
rect 3927 -16709 4000 -16705
rect 3927 -16757 3932 -16709
rect 3997 -16757 4000 -16709
rect 3927 -16762 4000 -16757
rect 2098 -17023 2123 -16952
rect 2521 -17023 2548 -16953
rect 2947 -17023 2972 -16950
rect 3372 -17023 3397 -16941
rect 3796 -17023 3821 -16914
rect 1534 -17074 4169 -17023
rect 1534 -17077 1826 -17074
rect 2098 -17083 2123 -17074
rect 2521 -17094 2548 -17074
rect 2947 -17081 2972 -17074
rect 3796 -17085 3821 -17074
<< via1 >>
rect 1892 0 1970 78
rect 1892 -523 1970 -445
rect 1892 -1046 1970 -968
rect 1892 -1569 1970 -1491
rect 1892 -2092 1970 -2014
rect 1892 -2615 1970 -2537
rect 1892 -3138 1970 -3060
rect 1892 -3661 1970 -3583
rect 1892 -4184 1970 -4106
rect 1892 -4707 1970 -4629
rect 1892 -5230 1970 -5152
rect 1892 -5753 1970 -5675
rect 1892 -6276 1970 -6198
rect 1892 -6799 1970 -6721
rect 1892 -7322 1970 -7244
rect 1892 -7845 1970 -7767
rect 1892 -8368 1970 -8290
rect 1892 -8891 1970 -8813
rect 1892 -9414 1970 -9336
rect 1892 -9937 1970 -9859
rect 1892 -10460 1970 -10382
rect 1892 -10983 1970 -10905
rect 1892 -11506 1970 -11428
rect 1892 -12029 1970 -11951
rect 1892 -12552 1970 -12474
rect 1892 -13075 1970 -12997
rect 1892 -13598 1970 -13520
rect 1892 -14121 1970 -14043
rect 1892 -14644 1970 -14566
rect 1892 -15167 1970 -15089
rect 1892 -15690 1970 -15612
rect 1956 -16208 2029 -16125
rect 2236 -16356 2301 -16308
rect 2658 -16350 2725 -16301
rect 3083 -16352 3148 -16304
rect 3511 -16356 3576 -16308
rect 3932 -16352 3997 -16304
rect 2218 -16599 2288 -16555
rect 2645 -16598 2712 -16549
rect 3067 -16596 3137 -16552
rect 3492 -16594 3562 -16550
rect 3918 -16594 3988 -16550
rect 2233 -16755 2298 -16707
rect 2656 -16755 2723 -16706
rect 3083 -16750 3148 -16702
rect 3506 -16752 3571 -16704
rect 3932 -16757 3997 -16709
rect 2215 -16995 2286 -16952
rect 2639 -16990 2710 -16947
rect 3063 -16995 3134 -16952
rect 3489 -16992 3560 -16949
rect 3915 -16990 3986 -16947
<< metal2 >>
rect 1887 78 1979 83
rect 1887 0 1892 78
rect 1970 0 1979 78
rect 1887 -9 1979 0
rect 1887 -445 1979 -440
rect 1887 -523 1892 -445
rect 1970 -523 1979 -445
rect 1887 -532 1979 -523
rect 1887 -968 1979 -963
rect 1887 -1046 1892 -968
rect 1970 -1046 1979 -968
rect 1887 -1055 1979 -1046
rect 1887 -1491 1979 -1486
rect 1887 -1569 1892 -1491
rect 1970 -1569 1979 -1491
rect 1887 -1578 1979 -1569
rect 1887 -2014 1979 -2009
rect 1887 -2092 1892 -2014
rect 1970 -2092 1979 -2014
rect 1887 -2101 1979 -2092
rect 1887 -2537 1979 -2532
rect 1887 -2615 1892 -2537
rect 1970 -2615 1979 -2537
rect 1887 -2624 1979 -2615
rect 1887 -3060 1979 -3055
rect 1887 -3138 1892 -3060
rect 1970 -3138 1979 -3060
rect 1887 -3147 1979 -3138
rect 1887 -3583 1979 -3578
rect 1887 -3661 1892 -3583
rect 1970 -3661 1979 -3583
rect 1887 -3670 1979 -3661
rect 1887 -4106 1979 -4101
rect 1887 -4184 1892 -4106
rect 1970 -4184 1979 -4106
rect 1887 -4193 1979 -4184
rect 1887 -4629 1979 -4624
rect 1887 -4707 1892 -4629
rect 1970 -4707 1979 -4629
rect 1887 -4716 1979 -4707
rect 1887 -5152 1979 -5147
rect 1887 -5230 1892 -5152
rect 1970 -5230 1979 -5152
rect 1887 -5239 1979 -5230
rect 1887 -5675 1979 -5670
rect 1887 -5753 1892 -5675
rect 1970 -5753 1979 -5675
rect 1887 -5762 1979 -5753
rect 1887 -6198 1979 -6193
rect 1887 -6276 1892 -6198
rect 1970 -6276 1979 -6198
rect 1887 -6285 1979 -6276
rect 1887 -6721 1979 -6716
rect 1887 -6799 1892 -6721
rect 1970 -6799 1979 -6721
rect 1887 -6808 1979 -6799
rect 1887 -7244 1979 -7239
rect 1887 -7322 1892 -7244
rect 1970 -7322 1979 -7244
rect 1887 -7331 1979 -7322
rect 1887 -7767 1979 -7762
rect 1887 -7845 1892 -7767
rect 1970 -7845 1979 -7767
rect 1887 -7854 1979 -7845
rect 1887 -8290 1979 -8285
rect 1887 -8368 1892 -8290
rect 1970 -8368 1979 -8290
rect 1887 -8377 1979 -8368
rect 1887 -8813 1979 -8808
rect 1887 -8891 1892 -8813
rect 1970 -8891 1979 -8813
rect 1887 -8900 1979 -8891
rect 1887 -9336 1979 -9331
rect 1887 -9414 1892 -9336
rect 1970 -9414 1979 -9336
rect 1887 -9423 1979 -9414
rect 1887 -9859 1979 -9854
rect 1887 -9937 1892 -9859
rect 1970 -9937 1979 -9859
rect 1887 -9946 1979 -9937
rect 1887 -10382 1979 -10377
rect 1887 -10460 1892 -10382
rect 1970 -10460 1979 -10382
rect 1887 -10469 1979 -10460
rect 1887 -10905 1979 -10900
rect 1887 -10983 1892 -10905
rect 1970 -10983 1979 -10905
rect 1887 -10992 1979 -10983
rect 1887 -11428 1979 -11423
rect 1887 -11506 1892 -11428
rect 1970 -11506 1979 -11428
rect 1887 -11515 1979 -11506
rect 1887 -11951 1979 -11946
rect 1887 -12029 1892 -11951
rect 1970 -12029 1979 -11951
rect 1887 -12038 1979 -12029
rect 1887 -12474 1979 -12469
rect 1887 -12552 1892 -12474
rect 1970 -12552 1979 -12474
rect 1887 -12561 1979 -12552
rect 1887 -12997 1979 -12992
rect 1887 -13075 1892 -12997
rect 1970 -13075 1979 -12997
rect 1887 -13084 1979 -13075
rect 1887 -13520 1979 -13515
rect 1887 -13598 1892 -13520
rect 1970 -13598 1979 -13520
rect 1887 -13607 1979 -13598
rect 1887 -14043 1979 -14038
rect 1887 -14121 1892 -14043
rect 1970 -14121 1979 -14043
rect 1887 -14130 1979 -14121
rect 1887 -14566 1979 -14561
rect 1887 -14644 1892 -14566
rect 1970 -14644 1979 -14566
rect 1887 -14653 1979 -14644
rect 1887 -15089 1979 -15084
rect 1887 -15167 1892 -15089
rect 1970 -15167 1979 -15089
rect 1887 -15176 1979 -15167
rect 1887 -15612 1979 -15607
rect 1887 -15690 1892 -15612
rect 1970 -15690 1979 -15612
rect 1887 -15699 1979 -15690
rect 1947 -16125 2039 -16116
rect 1947 -16208 1956 -16125
rect 2029 -16208 2039 -16125
rect 1947 -16217 2039 -16208
rect 2044 -16310 2165 -16247
rect 2230 -16306 2302 -16252
rect 2440 -16284 2593 -16236
rect 2230 -16308 2304 -16306
rect 2044 -16380 2121 -16310
rect 2230 -16317 2236 -16308
rect 2301 -16356 2304 -16308
rect 2440 -16350 2500 -16284
rect 2236 -16363 2304 -16356
rect 2439 -16361 2500 -16350
rect 2652 -16300 2724 -16236
rect 2903 -16259 3015 -16245
rect 2901 -16289 3015 -16259
rect 2652 -16301 2729 -16300
rect 2652 -16350 2658 -16301
rect 2725 -16350 2729 -16301
rect 2652 -16357 2729 -16350
rect 2653 -16358 2729 -16357
rect 2236 -16365 2270 -16363
rect 2046 -16621 2120 -16380
rect 2215 -16555 2290 -16551
rect 2215 -16599 2218 -16555
rect 2288 -16599 2290 -16555
rect 2215 -16603 2290 -16599
rect 2231 -16621 2281 -16603
rect 2046 -16680 2281 -16621
rect 2231 -16702 2281 -16680
rect 2439 -16634 2499 -16361
rect 2901 -16373 2973 -16289
rect 3087 -16301 3148 -16247
rect 3315 -16298 3441 -16250
rect 3080 -16304 3153 -16301
rect 3080 -16315 3083 -16304
rect 3148 -16352 3153 -16304
rect 3083 -16358 3153 -16352
rect 3315 -16366 3395 -16298
rect 3504 -16308 3579 -16245
rect 3737 -16250 3867 -16240
rect 3504 -16356 3511 -16308
rect 3576 -16356 3579 -16308
rect 3504 -16359 3579 -16356
rect 3506 -16361 3579 -16359
rect 3735 -16298 3867 -16250
rect 3735 -16364 3810 -16298
rect 3928 -16301 4000 -16252
rect 3928 -16304 4002 -16301
rect 3928 -16352 3932 -16304
rect 3997 -16352 4002 -16304
rect 3928 -16358 4002 -16352
rect 3928 -16359 4000 -16358
rect 2640 -16549 2716 -16545
rect 2640 -16598 2645 -16549
rect 2712 -16587 2716 -16549
rect 2712 -16598 2717 -16587
rect 2640 -16603 2717 -16598
rect 2656 -16634 2717 -16603
rect 2439 -16686 2717 -16634
rect 2901 -16613 2972 -16373
rect 3065 -16552 3140 -16547
rect 3065 -16596 3067 -16552
rect 3137 -16596 3140 -16552
rect 3065 -16599 3140 -16596
rect 3083 -16613 3139 -16599
rect 2901 -16669 3139 -16613
rect 2656 -16702 2717 -16686
rect 3083 -16700 3139 -16669
rect 3316 -16621 3393 -16366
rect 3490 -16550 3565 -16547
rect 3490 -16594 3492 -16550
rect 3562 -16594 3565 -16550
rect 3490 -16599 3565 -16594
rect 3504 -16621 3560 -16599
rect 3316 -16685 3560 -16621
rect 3504 -16700 3560 -16685
rect 3735 -16630 3803 -16364
rect 3916 -16550 3991 -16547
rect 3916 -16594 3918 -16550
rect 3988 -16594 3991 -16550
rect 3916 -16599 3991 -16594
rect 3929 -16630 3985 -16599
rect 3735 -16694 3985 -16630
rect 3078 -16702 3151 -16700
rect 2229 -16707 2302 -16702
rect 2229 -16755 2233 -16707
rect 2298 -16755 2302 -16707
rect 2229 -16759 2302 -16755
rect 2653 -16706 2729 -16702
rect 2653 -16755 2656 -16706
rect 2723 -16755 2729 -16706
rect 2653 -16760 2729 -16755
rect 3078 -16750 3083 -16702
rect 3148 -16750 3151 -16702
rect 3078 -16757 3151 -16750
rect 3502 -16704 3575 -16700
rect 3502 -16752 3506 -16704
rect 3571 -16752 3575 -16704
rect 3502 -16757 3575 -16752
rect 3927 -16705 3985 -16694
rect 3927 -16709 4000 -16705
rect 3927 -16757 3932 -16709
rect 3997 -16757 4000 -16709
rect 3927 -16762 4000 -16757
rect 2634 -16947 2719 -16933
rect 2212 -16952 2297 -16947
rect 2212 -16995 2215 -16952
rect 2286 -16995 2297 -16952
rect 2212 -17155 2297 -16995
rect 2634 -16990 2639 -16947
rect 2710 -16990 2719 -16947
rect 2634 -17141 2719 -16990
rect 3061 -16952 3146 -16947
rect 3061 -16995 3063 -16952
rect 3134 -16995 3146 -16952
rect 3061 -17155 3146 -16995
rect 3478 -16949 3563 -16942
rect 3478 -16992 3489 -16949
rect 3560 -16992 3563 -16949
rect 3478 -17150 3563 -16992
rect 3909 -16947 3994 -16942
rect 3909 -16990 3915 -16947
rect 3986 -16990 3994 -16947
rect 3909 -17150 3994 -16990
<< via2 >>
rect 1892 0 1970 78
rect 1892 -523 1970 -445
rect 1892 -1046 1970 -968
rect 1892 -1569 1970 -1491
rect 1892 -2092 1970 -2014
rect 1892 -2615 1970 -2537
rect 1892 -3138 1970 -3060
rect 1892 -3661 1970 -3583
rect 1892 -4184 1970 -4106
rect 1892 -4707 1970 -4629
rect 1892 -5230 1970 -5152
rect 1892 -5753 1970 -5675
rect 1892 -6276 1970 -6198
rect 1892 -6799 1970 -6721
rect 1892 -7322 1970 -7244
rect 1892 -7845 1970 -7767
rect 1892 -8368 1970 -8290
rect 1892 -8891 1970 -8813
rect 1892 -9414 1970 -9336
rect 1892 -9937 1970 -9859
rect 1892 -10460 1970 -10382
rect 1892 -10983 1970 -10905
rect 1892 -11506 1970 -11428
rect 1892 -12029 1970 -11951
rect 1892 -12552 1970 -12474
rect 1892 -13075 1970 -12997
rect 1892 -13598 1970 -13520
rect 1892 -14121 1970 -14043
rect 1892 -14644 1970 -14566
rect 1892 -15167 1970 -15089
rect 1892 -15690 1970 -15612
rect 1956 -16208 2029 -16125
<< metal3 >>
rect 1006 198 1477 515
rect 1006 146 3284 198
rect 1006 83 1477 146
rect 1006 78 1979 83
rect 1006 0 1892 78
rect 1970 0 1979 78
rect 1006 -9 1979 0
rect 1006 -440 1477 -9
rect 1006 -445 1979 -440
rect 1006 -523 1892 -445
rect 1970 -523 1979 -445
rect 1006 -532 1979 -523
rect 1006 -864 1477 -532
rect 1006 -916 3276 -864
rect 1006 -963 1477 -916
rect 1006 -968 1979 -963
rect 1006 -1046 1892 -968
rect 1970 -1046 1979 -968
rect 1006 -1055 1979 -1046
rect 1006 -1486 1477 -1055
rect 1006 -1491 1979 -1486
rect 1006 -1569 1892 -1491
rect 1970 -1569 1979 -1491
rect 1006 -1578 1979 -1569
rect 1006 -1906 1477 -1578
rect 1006 -1958 3288 -1906
rect 1006 -2009 1477 -1958
rect 1006 -2014 1979 -2009
rect 1006 -2092 1892 -2014
rect 1970 -2092 1979 -2014
rect 1006 -2101 1979 -2092
rect 1006 -2532 1477 -2101
rect 1006 -2537 1979 -2532
rect 1006 -2615 1892 -2537
rect 1970 -2615 1979 -2537
rect 1006 -2624 1979 -2615
rect 1006 -2956 1477 -2624
rect 1006 -3008 2920 -2956
rect 1006 -3055 1477 -3008
rect 1006 -3060 1979 -3055
rect 1006 -3138 1892 -3060
rect 1970 -3138 1979 -3060
rect 1006 -3147 1979 -3138
rect 1006 -3578 1477 -3147
rect 1006 -3583 1979 -3578
rect 1006 -3661 1892 -3583
rect 1970 -3661 1979 -3583
rect 1006 -3670 1979 -3661
rect 1006 -3994 1477 -3670
rect 1006 -4046 2956 -3994
rect 1006 -4101 1477 -4046
rect 1006 -4106 1979 -4101
rect 1006 -4184 1892 -4106
rect 1970 -4184 1979 -4106
rect 1006 -4193 1979 -4184
rect 1006 -4624 1477 -4193
rect 1006 -4629 1979 -4624
rect 1006 -4707 1892 -4629
rect 1970 -4707 1979 -4629
rect 1006 -4716 1979 -4707
rect 1006 -5044 1477 -4716
rect 1006 -5096 2908 -5044
rect 1006 -5147 1477 -5096
rect 1006 -5152 1979 -5147
rect 1006 -5230 1892 -5152
rect 1970 -5230 1979 -5152
rect 1006 -5239 1979 -5230
rect 1006 -5670 1477 -5239
rect 1006 -5675 1979 -5670
rect 1006 -5753 1892 -5675
rect 1970 -5753 1979 -5675
rect 1006 -5762 1979 -5753
rect 1006 -6086 1477 -5762
rect 1006 -6138 3256 -6086
rect 1006 -6193 1477 -6138
rect 1006 -6198 1979 -6193
rect 1006 -6276 1892 -6198
rect 1970 -6276 1979 -6198
rect 1006 -6285 1979 -6276
rect 1006 -6716 1477 -6285
rect 1006 -6721 1979 -6716
rect 1006 -6799 1892 -6721
rect 1970 -6799 1979 -6721
rect 1006 -6808 1979 -6799
rect 1006 -7136 1477 -6808
rect 1006 -7188 3264 -7136
rect 1006 -7239 1477 -7188
rect 1006 -7244 1979 -7239
rect 1006 -7322 1892 -7244
rect 1970 -7322 1979 -7244
rect 1006 -7331 1979 -7322
rect 1006 -7762 1477 -7331
rect 1006 -7767 1979 -7762
rect 1006 -7845 1892 -7767
rect 1970 -7845 1979 -7767
rect 1006 -7854 1979 -7845
rect 1006 -8186 1477 -7854
rect 1006 -8238 3264 -8186
rect 1006 -8285 1477 -8238
rect 1006 -8290 1979 -8285
rect 1006 -8368 1892 -8290
rect 1970 -8368 1979 -8290
rect 1006 -8377 1979 -8368
rect 1006 -8808 1477 -8377
rect 1006 -8813 1979 -8808
rect 1006 -8891 1892 -8813
rect 1970 -8891 1979 -8813
rect 1006 -8900 1979 -8891
rect 1006 -9216 1477 -8900
rect 1006 -9268 3288 -9216
rect 1006 -9331 1477 -9268
rect 1006 -9336 1979 -9331
rect 1006 -9414 1892 -9336
rect 1970 -9414 1979 -9336
rect 1006 -9423 1979 -9414
rect 1006 -9854 1477 -9423
rect 1006 -9859 1979 -9854
rect 1006 -9937 1892 -9859
rect 1970 -9937 1979 -9859
rect 1006 -9946 1979 -9937
rect 1006 -10262 1477 -9946
rect 1006 -10314 3288 -10262
rect 1006 -10377 1477 -10314
rect 1006 -10382 1979 -10377
rect 1006 -10460 1892 -10382
rect 1970 -10460 1979 -10382
rect 1006 -10469 1979 -10460
rect 1006 -10900 1477 -10469
rect 1006 -10905 1979 -10900
rect 1006 -10983 1892 -10905
rect 1970 -10983 1979 -10905
rect 1006 -10992 1979 -10983
rect 1006 -11324 1477 -10992
rect 1006 -11376 2948 -11324
rect 1006 -11423 1477 -11376
rect 1006 -11428 1979 -11423
rect 1006 -11506 1892 -11428
rect 1970 -11506 1979 -11428
rect 1006 -11515 1979 -11506
rect 1006 -11946 1477 -11515
rect 1006 -11951 1979 -11946
rect 1006 -12029 1892 -11951
rect 1970 -12029 1979 -11951
rect 1006 -12038 1979 -12029
rect 1006 -12357 1477 -12038
rect 1006 -12409 2900 -12357
rect 1006 -12469 1477 -12409
rect 1006 -12474 1979 -12469
rect 1006 -12552 1892 -12474
rect 1970 -12552 1979 -12474
rect 1006 -12561 1979 -12552
rect 1006 -12992 1477 -12561
rect 1006 -12997 1979 -12992
rect 1006 -13075 1892 -12997
rect 1970 -13075 1979 -12997
rect 1006 -13084 1979 -13075
rect 1006 -13403 1477 -13084
rect 1006 -13455 2888 -13403
rect 1006 -13515 1477 -13455
rect 1006 -13520 1979 -13515
rect 1006 -13598 1892 -13520
rect 1970 -13598 1979 -13520
rect 1006 -13607 1979 -13598
rect 1006 -14038 1477 -13607
rect 1006 -14043 1979 -14038
rect 1006 -14121 1892 -14043
rect 1970 -14121 1979 -14043
rect 1006 -14130 1979 -14121
rect 1006 -14453 1477 -14130
rect 1006 -14505 3260 -14453
rect 1006 -14561 1477 -14505
rect 1006 -14566 1979 -14561
rect 1006 -14644 1892 -14566
rect 1970 -14644 1979 -14566
rect 1006 -14653 1979 -14644
rect 1006 -15084 1477 -14653
rect 1006 -15089 1979 -15084
rect 1006 -15167 1892 -15089
rect 1970 -15167 1979 -15089
rect 1006 -15176 1979 -15167
rect 1006 -15499 1477 -15176
rect 1006 -15551 3260 -15499
rect 1006 -15607 1477 -15551
rect 1006 -15612 1979 -15607
rect 1006 -15690 1892 -15612
rect 1970 -15690 1979 -15612
rect 1006 -15699 1979 -15690
rect 1006 -16020 1477 -15699
rect 1006 -16072 2911 -16020
rect 1006 -16120 1477 -16072
rect 1947 -16120 2039 -16116
rect 1006 -16125 2039 -16120
rect 1006 -16208 1956 -16125
rect 2029 -16208 2039 -16125
rect 1006 -16212 2039 -16208
rect 1006 -17055 1477 -16212
rect 1947 -16217 2039 -16212
rect 2349 -17055 2426 -16451
rect 2772 -17055 2849 -16467
rect 3198 -17055 3275 -16465
rect 3619 -17055 3696 -16471
rect 4047 -17055 4124 -16476
rect 4157 -17055 4361 477
rect 1006 -17300 4415 -17055
use pbulk  pbulk_32 ~/Desktop/BENG207_Project/cochlea_sky130/mag/HW4_layout/3x8
timestamp 1639210801
transform 0 -1 2158 1 0 -16701
box -18 -18 119 75
use inv_customized_3  inv_customized_3_9
timestamp 1639205400
transform 0 -1 2552 1 0 -16515
box -85 128 180 481
use inv_customized_3  inv_customized_3_6
timestamp 1639205400
transform 0 -1 2550 1 0 -16916
box -85 128 180 481
use pbulk  pbulk_33
timestamp 1639210801
transform 0 -1 2594 1 0 -16701
box -18 -18 119 75
use inv_customized_3  inv_customized_3_8
timestamp 1639205400
transform 0 -1 2975 1 0 -16916
box -85 128 180 481
use inv_customized_3  inv_customized_3_7
timestamp 1639205400
transform 0 -1 2977 1 0 -16515
box -85 128 180 481
use pbulk  pbulk_34
timestamp 1639210801
transform 0 -1 3013 1 0 -16701
box -18 -18 119 75
use inv_customized_3  inv_customized_3_1
timestamp 1639205400
transform 0 -1 3402 1 0 -16515
box -85 128 180 481
use inv_customized_3  inv_customized_3_0
timestamp 1639205400
transform 0 -1 3400 1 0 -16916
box -85 128 180 481
use pbulk  pbulk_35
timestamp 1639210801
transform 0 -1 3442 1 0 -16709
box -18 -18 119 75
use inv_customized_3  inv_customized_3_3
timestamp 1639205400
transform 0 -1 3827 1 0 -16515
box -85 128 180 481
use inv_customized_3  inv_customized_3_2
timestamp 1639205400
transform 0 -1 3825 1 0 -16916
box -85 128 180 481
use pbulk  pbulk_36
timestamp 1639210801
transform 0 -1 3866 1 0 -16701
box -18 -18 119 75
use inv_customized_3  inv_customized_3_5
timestamp 1639205400
transform 0 -1 4252 1 0 -16515
box -85 128 180 481
use inv_customized_3  inv_customized_3_4
timestamp 1639205400
transform 0 -1 4250 1 0 -16916
box -85 128 180 481
use 0  0_159
timestamp 1639200303
transform -1 0 2330 0 1 -16321
box -89 43 336 566
use 0  0_143
timestamp 1639200303
transform 1 0 2508 0 1 -16321
box -89 43 336 566
use nbulk  nbulk_17
timestamp 1639219942
transform 1 0 2794 0 1 -16127
box -35 6 106 113
use 0  0_142
timestamp 1639200303
transform 1 0 2933 0 1 -16321
box -89 43 336 566
use 0  0_141
timestamp 1639200303
transform 1 0 3358 0 1 -16321
box -89 43 336 566
use 0  0_140
timestamp 1639200303
transform 1 0 3783 0 1 -16321
box -89 43 336 566
use inv_customized  inv_customized_16
timestamp 1639201766
transform 1 0 4309 0 1 -16324
box -194 128 180 481
use 0  0_158
timestamp 1639200303
transform -1 0 2330 0 1 -15798
box -89 43 336 566
use 0  0_139
timestamp 1639200303
transform 1 0 2508 0 1 -15798
box -89 43 336 566
use 0  0_138
timestamp 1639200303
transform 1 0 2933 0 1 -15798
box -89 43 336 566
use nbulk  nbulk_16
timestamp 1639219942
transform 1 0 3218 0 1 -15599
box -35 6 106 113
use pbulk  pbulk_31
timestamp 1639210801
transform 1 0 3094 0 1 -15889
box -18 -18 119 75
use 0  0_137
timestamp 1639200303
transform 1 0 3358 0 1 -15798
box -89 43 336 566
use 0  0_136
timestamp 1639200303
transform -1 0 4030 0 1 -15798
box -89 43 336 566
use inv_customized  inv_customized_17
timestamp 1639201766
transform 1 0 4309 0 1 -15801
box -194 128 180 481
use 0  0_157
timestamp 1639200303
transform -1 0 2330 0 1 -15275
box -89 43 336 566
use 0  0_133
timestamp 1639200303
transform 1 0 2508 0 1 -15275
box -89 43 336 566
use 0  0_134
timestamp 1639200303
transform 1 0 2933 0 1 -15275
box -89 43 336 566
use 0  0_135
timestamp 1639200303
transform -1 0 3605 0 1 -15275
box -89 43 336 566
use pbulk  pbulk_30
timestamp 1639210801
transform 1 0 3654 0 1 -15377
box -18 -18 119 75
use 0  0_132
timestamp 1639200303
transform -1 0 4030 0 1 -15275
box -89 43 336 566
use inv_customized  inv_customized_18
timestamp 1639201766
transform 1 0 4309 0 1 -15278
box -194 128 180 481
use 0  0_156
timestamp 1639200303
transform -1 0 2330 0 1 -14752
box -89 43 336 566
use 0  0_130
timestamp 1639200303
transform 1 0 2508 0 1 -14752
box -89 43 336 566
use 0  0_129
timestamp 1639200303
transform 1 0 2933 0 1 -14752
box -89 43 336 566
use nbulk  nbulk_15
timestamp 1639219942
transform 1 0 3230 0 1 -14545
box -35 6 106 113
use pbulk  pbulk_29
timestamp 1639210801
transform 1 0 3240 0 1 -14853
box -18 -18 119 75
use 0  0_131
timestamp 1639200303
transform -1 0 3605 0 1 -14752
box -89 43 336 566
use 0  0_128
timestamp 1639200303
transform 1 0 3783 0 1 -14752
box -89 43 336 566
use inv_customized  inv_customized_19
timestamp 1639201766
transform 1 0 4309 0 1 -14755
box -194 128 180 481
use 0  0_155
timestamp 1639200303
transform -1 0 2330 0 1 -14229
box -89 43 336 566
use 0  0_127
timestamp 1639200303
transform 1 0 2508 0 1 -14229
box -89 43 336 566
use 0  0_126
timestamp 1639200303
transform -1 0 3180 0 1 -14229
box -89 43 336 566
use pbulk  pbulk_28
timestamp 1639210801
transform 1 0 3166 0 1 -14330
box -18 -18 119 75
use 0  0_125
timestamp 1639200303
transform -1 0 3605 0 1 -14229
box -89 43 336 566
use 0  0_124
timestamp 1639200303
transform 1 0 3783 0 1 -14229
box -89 43 336 566
use inv_customized  inv_customized_20
timestamp 1639201766
transform 1 0 4309 0 1 -14232
box -194 128 180 481
use 0  0_154
timestamp 1639200303
transform -1 0 2330 0 1 -13706
box -89 43 336 566
use 0  0_121
timestamp 1639200303
transform 1 0 2508 0 1 -13706
box -89 43 336 566
use nbulk  nbulk_14
timestamp 1639219942
transform 1 0 2810 0 1 -13495
box -35 6 106 113
use pbulk  pbulk_27
timestamp 1639210801
transform 1 0 2811 0 1 -13806
box -18 -18 119 75
use 0  0_122
timestamp 1639200303
transform -1 0 3180 0 1 -13706
box -89 43 336 566
use 0  0_123
timestamp 1639200303
transform -1 0 3605 0 1 -13706
box -89 43 336 566
use 0  0_120
timestamp 1639200303
transform -1 0 4030 0 1 -13706
box -89 43 336 566
use inv_customized  inv_customized_21
timestamp 1639201766
transform 1 0 4309 0 1 -13709
box -194 128 180 481
use 0  0_153
timestamp 1639200303
transform -1 0 2330 0 1 -13183
box -89 43 336 566
use 0  0_119
timestamp 1639200303
transform 1 0 2508 0 1 -13183
box -89 43 336 566
use pbulk  pbulk_26
timestamp 1639210801
transform 1 0 2804 0 1 -13280
box -18 -18 119 75
use 0  0_118
timestamp 1639200303
transform -1 0 3180 0 1 -13183
box -89 43 336 566
use 0  0_117
timestamp 1639200303
transform 1 0 3358 0 1 -13183
box -89 43 336 566
use 0  0_116
timestamp 1639200303
transform -1 0 4030 0 1 -13183
box -89 43 336 566
use inv_customized  inv_customized_22
timestamp 1639201766
transform 1 0 4309 0 1 -13186
box -194 128 180 481
use 0  0_152
timestamp 1639200303
transform -1 0 2330 0 1 -12660
box -89 43 336 566
use 0  0_113
timestamp 1639200303
transform 1 0 2508 0 1 -12660
box -89 43 336 566
use nbulk  nbulk_13
timestamp 1639219942
transform 1 0 2808 0 1 -12453
box -35 6 106 113
use pbulk  pbulk_25
timestamp 1639210801
transform 1 0 2809 0 1 -12766
box -18 -18 119 75
use 0  0_114
timestamp 1639200303
transform -1 0 3180 0 1 -12660
box -89 43 336 566
use 0  0_115
timestamp 1639200303
transform 1 0 3358 0 1 -12660
box -89 43 336 566
use 0  0_112
timestamp 1639200303
transform 1 0 3783 0 1 -12660
box -89 43 336 566
use inv_customized  inv_customized_23
timestamp 1639201766
transform 1 0 4309 0 1 -12663
box -194 128 180 481
use 0  0_151
timestamp 1639200303
transform -1 0 2330 0 1 -12137
box -89 43 336 566
use 0  0_111
timestamp 1639200303
transform -1 0 2755 0 1 -12137
box -89 43 336 566
use pbulk  pbulk_24
timestamp 1639210801
transform 1 0 2806 0 1 -12238
box -18 -18 119 75
use 0  0_110
timestamp 1639200303
transform -1 0 3180 0 1 -12137
box -89 43 336 566
use 0  0_109
timestamp 1639200303
transform 1 0 3358 0 1 -12137
box -89 43 336 566
use 0  0_108
timestamp 1639200303
transform 1 0 3783 0 1 -12137
box -89 43 336 566
use inv_customized  inv_customized_25
timestamp 1639201766
transform 1 0 4309 0 1 -12140
box -194 128 180 481
use pbulk  pbulk_23
timestamp 1639210801
transform 1 0 2395 0 1 -11714
box -18 -18 119 75
use 0  0_150
timestamp 1639200303
transform -1 0 2330 0 1 -11614
box -89 43 336 566
use 0  0_107
timestamp 1639200303
transform -1 0 2755 0 1 -11614
box -89 43 336 566
use nbulk  nbulk_12
timestamp 1639219942
transform 1 0 2840 0 1 -11411
box -35 6 106 113
use 0  0_106
timestamp 1639200303
transform -1 0 3180 0 1 -11614
box -89 43 336 566
use 0  0_105
timestamp 1639200303
transform 1 0 3358 0 1 -11614
box -89 43 336 566
use 0  0_104
timestamp 1639200303
transform -1 0 4030 0 1 -11614
box -89 43 336 566
use inv_customized  inv_customized_24
timestamp 1639201766
transform 1 0 4309 0 1 -11617
box -194 128 180 481
use 0  0_149
timestamp 1639200303
transform -1 0 2330 0 1 -11091
box -89 43 336 566
use 0  0_103
timestamp 1639200303
transform -1 0 2755 0 1 -11091
box -89 43 336 566
use 0  0_102
timestamp 1639200303
transform -1 0 3180 0 1 -11091
box -89 43 336 566
use 0  0_101
timestamp 1639200303
transform -1 0 3605 0 1 -11091
box -89 43 336 566
use pbulk  pbulk_22
timestamp 1639210801
transform 1 0 3659 0 1 -11193
box -18 -18 119 75
use 0  0_100
timestamp 1639200303
transform -1 0 4030 0 1 -11091
box -89 43 336 566
use inv_customized  inv_customized_27
timestamp 1639201766
transform 1 0 4309 0 1 -11094
box -194 128 180 481
use 0  0_148
timestamp 1639200303
transform -1 0 2330 0 1 -10568
box -89 43 336 566
use 0  0_97
timestamp 1639200303
transform -1 0 2755 0 1 -10568
box -89 43 336 566
use 0  0_98
timestamp 1639200303
transform -1 0 3180 0 1 -10568
box -89 43 336 566
use nbulk  nbulk_11
timestamp 1639219942
transform 1 0 3268 0 1 -10357
box -35 6 106 113
use pbulk  pbulk_21
timestamp 1639210801
transform 1 0 3249 0 1 -10667
box -18 -18 119 75
use 0  0_99
timestamp 1639200303
transform -1 0 3605 0 1 -10568
box -89 43 336 566
use 0  0_96
timestamp 1639200303
transform 1 0 3783 0 1 -10568
box -89 43 336 566
use inv_customized  inv_customized_26
timestamp 1639201766
transform 1 0 4309 0 1 -10571
box -194 128 180 481
use 0  0_147
timestamp 1639200303
transform -1 0 2330 0 1 -10045
box -89 43 336 566
use 0  0_95
timestamp 1639200303
transform -1 0 2755 0 1 -10045
box -89 43 336 566
use 0  0_94
timestamp 1639200303
transform 1 0 2933 0 1 -10045
box -89 43 336 566
use pbulk  pbulk_20
timestamp 1639210801
transform 1 0 3278 0 1 -10146
box -18 -18 119 75
use 0  0_93
timestamp 1639200303
transform -1 0 3605 0 1 -10045
box -89 43 336 566
use 0  0_92
timestamp 1639200303
transform 1 0 3783 0 1 -10045
box -89 43 336 566
use inv_customized  inv_customized_29
timestamp 1639201766
transform 1 0 4309 0 1 -10048
box -194 128 180 481
use 0  0_146
timestamp 1639200303
transform -1 0 2330 0 1 -9522
box -89 43 336 566
use 0  0_91
timestamp 1639200303
transform -1 0 2755 0 1 -9522
box -89 43 336 566
use 0  0_90
timestamp 1639200303
transform 1 0 2933 0 1 -9522
box -89 43 336 566
use nbulk  nbulk_10
timestamp 1639219942
transform 1 0 3240 0 1 -9313
box -35 6 106 113
use pbulk  pbulk_19
timestamp 1639210801
transform 1 0 3228 0 1 -9622
box -18 -18 119 75
use 0  0_89
timestamp 1639200303
transform -1 0 3605 0 1 -9522
box -89 43 336 566
use 0  0_88
timestamp 1639200303
transform -1 0 4030 0 1 -9522
box -89 43 336 566
use inv_customized  inv_customized_28
timestamp 1639201766
transform 1 0 4309 0 1 -9525
box -194 128 180 481
use 0  0_145
timestamp 1639200303
transform -1 0 2330 0 1 -8999
box -89 43 336 566
use 0  0_87
timestamp 1639200303
transform -1 0 2755 0 1 -8999
box -89 43 336 566
use 0  0_86
timestamp 1639200303
transform 1 0 2933 0 1 -8999
box -89 43 336 566
use pbulk  pbulk_18
timestamp 1639210801
transform 1 0 3218 0 1 -9101
box -18 -18 119 75
use 0  0_85
timestamp 1639200303
transform 1 0 3358 0 1 -8999
box -89 43 336 566
use 0  0_84
timestamp 1639200303
transform -1 0 4030 0 1 -8999
box -89 43 336 566
use inv_customized  inv_customized_30
timestamp 1639201766
transform 1 0 4309 0 1 -9002
box -194 128 180 481
use 0  0_144
timestamp 1639200303
transform -1 0 2330 0 1 -8476
box -89 43 336 566
use 0  0_83
timestamp 1639200303
transform -1 0 2755 0 1 -8476
box -89 43 336 566
use 0  0_82
timestamp 1639200303
transform 1 0 2933 0 1 -8476
box -89 43 336 566
use nbulk  nbulk_9
timestamp 1639219942
transform 1 0 3210 0 1 -8281
box -35 6 106 113
use 0  0_81
timestamp 1639200303
transform 1 0 3358 0 1 -8476
box -89 43 336 566
use pbulk  pbulk_17
timestamp 1639210801
transform 1 0 3657 0 1 -8575
box -18 -18 119 75
use 0  0_80
timestamp 1639200303
transform 1 0 3783 0 1 -8476
box -89 43 336 566
use inv_customized  inv_customized_31
timestamp 1639201766
transform 1 0 4309 0 1 -8479
box -194 128 180 481
use pbulk  pbulk_16
timestamp 1639210801
transform 1 0 2422 0 1 -8054
box -18 -18 119 75
use 0  0_79
timestamp 1639200303
transform 1 0 2083 0 1 -7953
box -89 43 336 566
use 0  0_63
timestamp 1639200303
transform -1 0 2755 0 1 -7953
box -89 43 336 566
use 0  0_55
timestamp 1639200303
transform 1 0 2933 0 1 -7953
box -89 43 336 566
use 0  0_54
timestamp 1639200303
transform 1 0 3358 0 1 -7953
box -89 43 336 566
use 0  0_53
timestamp 1639200303
transform 1 0 3783 0 1 -7953
box -89 43 336 566
use inv_customized  inv_customized_15
timestamp 1639201766
transform 1 0 4309 0 1 -7956
box -194 128 180 481
use pbulk  pbulk_15
timestamp 1639210801
transform 1 0 2360 0 1 -7530
box -18 -18 119 75
use 0  0_78
timestamp 1639200303
transform 1 0 2083 0 1 -7430
box -89 43 336 566
use 0  0_62
timestamp 1639200303
transform -1 0 2755 0 1 -7430
box -89 43 336 566
use 0  0_50
timestamp 1639200303
transform 1 0 2933 0 1 -7430
box -89 43 336 566
use nbulk  nbulk_8
timestamp 1639219942
transform 1 0 3212 0 1 -7237
box -35 6 106 113
use 0  0_52
timestamp 1639200303
transform 1 0 3358 0 1 -7430
box -89 43 336 566
use 0  0_51
timestamp 1639200303
transform -1 0 4030 0 1 -7430
box -89 43 336 566
use inv_customized  inv_customized_8
timestamp 1639201766
transform 1 0 4309 0 1 -7433
box -194 128 180 481
use 0  0_77
timestamp 1639200303
transform 1 0 2083 0 1 -6907
box -89 43 336 566
use 0  0_61
timestamp 1639200303
transform -1 0 2755 0 1 -6907
box -89 43 336 566
use 0  0_47
timestamp 1639200303
transform 1 0 2933 0 1 -6907
box -89 43 336 566
use pbulk  pbulk_14
timestamp 1639210801
transform 1 0 3205 0 1 -7006
box -18 -18 119 75
use 0  0_49
timestamp 1639200303
transform -1 0 3605 0 1 -6907
box -89 43 336 566
use 0  0_48
timestamp 1639200303
transform -1 0 4030 0 1 -6907
box -89 43 336 566
use inv_customized  inv_customized_9
timestamp 1639201766
transform 1 0 4309 0 1 -6910
box -194 128 180 481
use 0  0_76
timestamp 1639200303
transform 1 0 2083 0 1 -6384
box -89 43 336 566
use 0  0_60
timestamp 1639200303
transform -1 0 2755 0 1 -6384
box -89 43 336 566
use 0  0_44
timestamp 1639200303
transform 1 0 2933 0 1 -6384
box -89 43 336 566
use nbulk  nbulk_7
timestamp 1639219942
transform 1 0 3234 0 1 -6177
box -35 6 106 113
use pbulk  pbulk_13
timestamp 1639210801
transform 1 0 3230 0 1 -6480
box -18 -18 119 75
use 0  0_46
timestamp 1639200303
transform -1 0 3605 0 1 -6384
box -89 43 336 566
use 0  0_45
timestamp 1639200303
transform 1 0 3783 0 1 -6384
box -89 43 336 566
use inv_customized  inv_customized_10
timestamp 1639201766
transform 1 0 4309 0 1 -6387
box -194 128 180 481
use 0  0_75
timestamp 1639200303
transform 1 0 2083 0 1 -5861
box -89 43 336 566
use 0  0_59
timestamp 1639200303
transform -1 0 2755 0 1 -5861
box -89 43 336 566
use 0  0_41
timestamp 1639200303
transform -1 0 3180 0 1 -5861
box -89 43 336 566
use pbulk  pbulk_12
timestamp 1639210801
transform 1 0 3223 0 1 -5959
box -18 -18 119 75
use 0  0_43
timestamp 1639200303
transform -1 0 3605 0 1 -5861
box -89 43 336 566
use 0  0_42
timestamp 1639200303
transform 1 0 3783 0 1 -5861
box -89 43 336 566
use inv_customized  inv_customized_11
timestamp 1639201766
transform 1 0 4309 0 1 -5864
box -194 128 180 481
use 0  0_74
timestamp 1639200303
transform 1 0 2083 0 1 -5338
box -89 43 336 566
use 0  0_58
timestamp 1639200303
transform -1 0 2755 0 1 -5338
box -89 43 336 566
use nbulk  nbulk_6
timestamp 1639219942
transform 1 0 2844 0 1 -5141
box -35 6 106 113
use pbulk  pbulk_11
timestamp 1639210801
transform 1 0 2846 0 1 -5441
box -18 -18 119 75
use 0  0_38
timestamp 1639200303
transform -1 0 3180 0 1 -5338
box -89 43 336 566
use 0  0_40
timestamp 1639200303
transform -1 0 3605 0 1 -5338
box -89 43 336 566
use 0  0_39
timestamp 1639200303
transform -1 0 4030 0 1 -5338
box -89 43 336 566
use inv_customized  inv_customized_12
timestamp 1639201766
transform 1 0 4309 0 1 -5341
box -194 128 180 481
use 0  0_73
timestamp 1639200303
transform 1 0 2083 0 1 -4815
box -89 43 336 566
use 0  0_57
timestamp 1639200303
transform -1 0 2755 0 1 -4815
box -89 43 336 566
use pbulk  pbulk_10
timestamp 1639210801
transform 1 0 2844 0 1 -4917
box -18 -18 119 75
use 0  0_35
timestamp 1639200303
transform -1 0 3180 0 1 -4815
box -89 43 336 566
use 0  0_37
timestamp 1639200303
transform 1 0 3358 0 1 -4815
box -89 43 336 566
use 0  0_36
timestamp 1639200303
transform -1 0 4030 0 1 -4815
box -89 43 336 566
use inv_customized  inv_customized_13
timestamp 1639201766
transform 1 0 4309 0 1 -4818
box -194 128 180 481
use 0  0_72
timestamp 1639200303
transform 1 0 2083 0 1 -4292
box -89 43 336 566
use 0  0_56
timestamp 1639200303
transform -1 0 2755 0 1 -4292
box -89 43 336 566
use nbulk  nbulk_5
timestamp 1639219942
transform 1 0 2850 0 1 -4089
box -35 6 106 113
use pbulk  pbulk_9
timestamp 1639210801
transform 1 0 2839 0 1 -4391
box -18 -18 119 75
use 0  0_32
timestamp 1639200303
transform -1 0 3180 0 1 -4292
box -89 43 336 566
use 0  0_34
timestamp 1639200303
transform 1 0 3358 0 1 -4292
box -89 43 336 566
use 0  0_33
timestamp 1639200303
transform 1 0 3783 0 1 -4292
box -89 43 336 566
use inv_customized  inv_customized_14
timestamp 1639201766
transform 1 0 4309 0 1 -4295
box -194 128 180 481
use 0  0_71
timestamp 1639200303
transform 1 0 2083 0 1 -3769
box -89 43 336 566
use 0  0_31
timestamp 1639200303
transform 1 0 2508 0 1 -3769
box -89 43 336 566
use pbulk  pbulk_8
timestamp 1639210801
transform 1 0 2841 0 1 -3870
box -18 -18 119 75
use 0  0_23
timestamp 1639200303
transform -1 0 3180 0 1 -3769
box -89 43 336 566
use 0  0_18
timestamp 1639200303
transform 1 0 3358 0 1 -3769
box -89 43 336 566
use 0  0_19
timestamp 1639200303
transform 1 0 3783 0 1 -3769
box -89 43 336 566
use inv_customized  inv_customized_7
timestamp 1639201766
transform 1 0 4309 0 1 -3772
box -194 128 180 481
use 0  0_70
timestamp 1639200303
transform 1 0 2083 0 1 -3246
box -89 43 336 566
use 0  0_30
timestamp 1639200303
transform 1 0 2508 0 1 -3246
box -89 43 336 566
use nbulk  nbulk_4
timestamp 1639219942
transform 1 0 2814 0 1 -3041
box -35 6 106 113
use pbulk  pbulk_7
timestamp 1639210801
transform 1 0 2799 0 1 -3346
box -18 -18 119 75
use 0  0_22
timestamp 1639200303
transform -1 0 3180 0 1 -3246
box -89 43 336 566
use 0  0_16
timestamp 1639200303
transform 1 0 3358 0 1 -3246
box -89 43 336 566
use 0  0_17
timestamp 1639200303
transform -1 0 4030 0 1 -3246
box -89 43 336 566
use inv_customized  inv_customized_6
timestamp 1639201766
transform 1 0 4309 0 1 -3249
box -194 128 180 481
use 0  0_69
timestamp 1639200303
transform 1 0 2083 0 1 -2723
box -89 43 336 566
use 0  0_29
timestamp 1639200303
transform 1 0 2508 0 1 -2723
box -89 43 336 566
use pbulk  pbulk_6
timestamp 1639210801
transform 1 0 2809 0 1 -2822
box -18 -18 119 75
use 0  0_21
timestamp 1639200303
transform -1 0 3180 0 1 -2723
box -89 43 336 566
use 0  0_15
timestamp 1639200303
transform -1 0 3605 0 1 -2723
box -89 43 336 566
use 0  0_14
timestamp 1639200303
transform -1 0 4030 0 1 -2723
box -89 43 336 566
use inv_customized  inv_customized_5
timestamp 1639201766
transform 1 0 4309 0 1 -2726
box -194 128 180 481
use 0  0_68
timestamp 1639200303
transform 1 0 2083 0 1 -2200
box -89 43 336 566
use 0  0_28
timestamp 1639200303
transform 1 0 2508 0 1 -2200
box -89 43 336 566
use pbulk  pbulk_5
timestamp 1639210801
transform 1 0 2796 0 1 -2299
box -18 -18 119 75
use 0  0_20
timestamp 1639200303
transform -1 0 3180 0 1 -2200
box -89 43 336 566
use nbulk  nbulk_3
timestamp 1639219942
transform 1 0 3266 0 1 -1993
box -35 6 106 113
use 0  0_12
timestamp 1639200303
transform -1 0 3605 0 1 -2200
box -89 43 336 566
use 0  0_13
timestamp 1639200303
transform 1 0 3783 0 1 -2200
box -89 43 336 566
use inv_customized  inv_customized_4
timestamp 1639201766
transform 1 0 4309 0 1 -2203
box -194 128 180 481
use 0  0_67
timestamp 1639200303
transform 1 0 2083 0 1 -1677
box -89 43 336 566
use 0  0_27
timestamp 1639200303
transform 1 0 2508 0 1 -1677
box -89 43 336 566
use pbulk  pbulk_4
timestamp 1639210801
transform 1 0 2789 0 1 -1773
box -18 -18 119 75
use 0  0_11
timestamp 1639200303
transform 1 0 2933 0 1 -1677
box -89 43 336 566
use 0  0_2
timestamp 1639200303
transform -1 0 3605 0 1 -1677
box -89 43 336 566
use 0  0_7
timestamp 1639200303
transform 1 0 3783 0 1 -1677
box -89 43 336 566
use inv_customized  inv_customized_3
timestamp 1639201766
transform 1 0 4309 0 1 -1680
box -194 128 180 481
use 0  0_66
timestamp 1639200303
transform 1 0 2083 0 1 -1154
box -89 43 336 566
use 0  0_26
timestamp 1639200303
transform 1 0 2508 0 1 -1154
box -89 43 336 566
use pbulk  pbulk_3
timestamp 1639210801
transform 1 0 2767 0 1 -1254
box -18 -18 119 75
use 0  0_10
timestamp 1639200303
transform 1 0 2933 0 1 -1154
box -89 43 336 566
use nbulk  nbulk_1
timestamp 1639219942
transform 1 0 3222 0 1 -949
box -35 6 106 113
use 0  0_4
timestamp 1639200303
transform -1 0 3605 0 1 -1154
box -89 43 336 566
use 0  0_6
timestamp 1639200303
transform -1 0 4030 0 1 -1154
box -89 43 336 566
use inv_customized  inv_customized_2
timestamp 1639201766
transform 1 0 4309 0 1 -1157
box -194 128 180 481
use 0  0_65
timestamp 1639200303
transform 1 0 2083 0 1 -631
box -89 43 336 566
use 0  0_25
timestamp 1639200303
transform 1 0 2508 0 1 -631
box -89 43 336 566
use pbulk  pbulk_2
timestamp 1639210801
transform 1 0 2757 0 1 -730
box -18 -18 119 75
use 0  0_9
timestamp 1639200303
transform 1 0 2933 0 1 -631
box -89 43 336 566
use 0  0_3
timestamp 1639200303
transform 1 0 3358 0 1 -631
box -89 43 336 566
use 0  0_5
timestamp 1639200303
transform -1 0 4030 0 1 -631
box -89 43 336 566
use inv_customized  inv_customized_1
timestamp 1639201766
transform 1 0 4309 0 1 -634
box -194 128 180 481
use 0  0_64
timestamp 1639200303
transform 1 0 2083 0 1 -108
box -89 43 336 566
use 0  0_24
timestamp 1639200303
transform 1 0 2508 0 1 -108
box -89 43 336 566
use pbulk  pbulk_1
timestamp 1639210801
transform 1 0 2779 0 1 -202
box -18 -18 119 75
use 0  0_8
timestamp 1639200303
transform 1 0 2933 0 1 -108
box -89 43 336 566
use nbulk  nbulk_0
timestamp 1639219942
transform 1 0 3186 0 1 109
box -35 6 106 113
use 0  0_0
timestamp 1639200303
transform 1 0 3358 0 1 -108
box -89 43 336 566
use 0  0_1
timestamp 1639200303
transform 1 0 3783 0 1 -108
box -89 43 336 566
use inv_customized  inv_customized_0
timestamp 1639201766
transform 1 0 4309 0 1 -111
box -194 128 180 481
use pbulk  pbulk_0
timestamp 1639210801
transform 1 0 2777 0 1 319
box -18 -18 119 75
<< labels >>
rlabel metal1 1996 -191 1996 -191 7 W1
port 1 w
rlabel metal1 1996 -714 1996 -714 7 W1
port 1 w
rlabel metal1 1996 -1237 1996 -1237 7 W1
port 1 w
rlabel metal1 1996 -1760 1996 -1760 7 W1
port 1 w
rlabel metal1 1996 -2283 1996 -2283 7 W1
port 1 w
rlabel metal1 1996 -2806 1996 -2806 7 W1
port 1 w
rlabel metal1 1996 -3329 1996 -3329 7 W1
port 1 w
rlabel metal1 1996 -3852 1996 -3852 7 W1
port 1 w
rlabel metal1 1996 -4375 1996 -4375 7 W1
port 1 w
rlabel metal1 1996 -4898 1996 -4898 7 W1
port 1 w
rlabel metal1 1996 -5421 1996 -5421 7 W1
port 1 w
rlabel metal1 1996 -5944 1996 -5944 7 W1
port 1 w
rlabel metal1 1996 -6467 1996 -6467 7 W1
port 1 w
rlabel metal1 1996 -6990 1996 -6990 7 W1
port 1 w
rlabel metal1 1996 -7513 1996 -7513 7 W1
port 1 w
rlabel metal1 1996 -8036 1996 -8036 7 W1
port 1 w
rlabel metal1 1996 -8559 1996 -8559 7 W1
port 1 w
rlabel metal1 1996 -9082 1996 -9082 7 W1
port 1 w
rlabel metal1 1996 -9605 1996 -9605 7 W1
port 1 w
rlabel metal1 1996 -10128 1996 -10128 7 W1
port 1 w
rlabel metal1 1996 -10651 1996 -10651 7 W1
port 1 w
rlabel metal1 1996 -11174 1996 -11174 7 W1
port 1 w
rlabel metal1 1996 -11697 1996 -11697 7 W1
port 1 w
rlabel metal1 1996 -12220 1996 -12220 7 W1
port 1 w
rlabel metal1 1996 -12743 1996 -12743 7 W1
port 1 w
rlabel metal1 1996 -13266 1996 -13266 7 W1
port 1 w
rlabel metal1 1996 -13789 1996 -13789 7 W1
port 1 w
rlabel metal1 1996 -14312 1996 -14312 7 W1
port 1 w
rlabel metal1 1996 -14835 1996 -14835 7 W1
port 1 w
rlabel metal1 1996 -15358 1996 -15358 7 W1
port 1 w
rlabel metal1 1996 -15881 1996 -15881 7 W1
port 1 w
rlabel metal1 1995 -475 1995 -475 7 W3
port 3 w
rlabel metal1 1995 -998 1995 -998 7 W3
port 3 w
rlabel metal1 1995 -1521 1995 -1521 7 W3
port 3 w
rlabel metal1 1995 -2044 1995 -2044 7 W3
port 3 w
rlabel metal1 1995 -2567 1995 -2567 7 W3
port 3 w
rlabel metal1 1995 -3090 1995 -3090 7 W3
port 3 w
rlabel metal1 1995 -3613 1995 -3613 7 W3
port 3 w
rlabel metal1 1995 -4136 1995 -4136 7 W3
port 3 w
rlabel metal1 1995 -4659 1995 -4659 7 W3
port 3 w
rlabel metal1 1995 -5182 1995 -5182 7 W3
port 3 w
rlabel metal1 1995 -5705 1995 -5705 7 W3
port 3 w
rlabel metal1 1995 -6228 1995 -6228 7 W3
port 3 w
rlabel metal1 1995 -6751 1995 -6751 7 W3
port 3 w
rlabel metal1 1995 -7274 1995 -7274 7 W3
port 3 w
rlabel metal1 1995 -7797 1995 -7797 7 W3
port 3 w
rlabel metal1 1995 -8320 1995 -8320 7 W3
port 3 w
rlabel metal1 1995 -8843 1995 -8843 7 W3
port 3 w
rlabel metal1 1995 -9366 1995 -9366 7 W3
port 3 w
rlabel metal1 1995 -9889 1995 -9889 7 W3
port 3 w
rlabel metal1 1995 -10412 1995 -10412 7 W3
port 3 w
rlabel metal1 1995 -10935 1995 -10935 7 W3
port 3 w
rlabel metal1 1995 -11458 1995 -11458 7 W3
port 3 w
rlabel metal1 1995 -11981 1995 -11981 7 W3
port 3 w
rlabel metal1 1995 -12504 1995 -12504 7 W3
port 3 w
rlabel metal1 1995 -13027 1995 -13027 7 W3
port 3 w
rlabel metal1 1995 -13550 1995 -13550 7 W3
port 3 w
rlabel metal1 1995 -14073 1995 -14073 7 W3
port 3 w
rlabel metal1 1995 -14596 1995 -14596 7 W3
port 3 w
rlabel metal1 1995 -15119 1995 -15119 7 W3
port 3 w
rlabel metal1 1995 -15642 1995 -15642 7 W3
port 3 w
rlabel space 4472 -16045 4472 -16045 1 sel0
rlabel space 4477 -15523 4477 -15523 1 sel1
rlabel space 4483 -14998 4483 -14998 1 sel2
rlabel space 4479 -14475 4479 -14475 1 sel3
rlabel space 4477 -13951 4477 -13951 1 sel4
rlabel space 4475 -13426 4475 -13426 1 sel5
rlabel space 4480 -12900 4480 -12900 1 sel6
rlabel space 4480 -12370 4480 -12370 1 sel7
rlabel space 4483 -11864 4483 -11864 1 sel8
rlabel space 4482 -11332 4482 -11332 1 sel9
rlabel space 4484 -10812 4484 -10812 7 sel10
rlabel space 4483 -10289 4483 -10289 1 sel11
rlabel space 4480 -9765 4480 -9765 1 sel12
rlabel space 4479 -9240 4479 -9240 1 sel13
rlabel space 4482 -8724 4482 -8724 1 sel14
rlabel space 4478 -8200 4478 -8200 1 sel15
rlabel space 4483 -7673 4483 -7673 1 sel16
rlabel space 4483 -7149 4483 -7149 1 sel17
rlabel space 4486 -6627 4486 -6627 7 sel18
rlabel space 4485 -6105 4485 -6105 7 sel19
rlabel space 4487 -5582 4487 -5582 7 sel20
rlabel space 4485 -5056 4485 -5056 7 sel21
rlabel space 4483 -4538 4483 -4538 1 sel22
rlabel space 4482 -4013 4482 -4013 1 sel23
rlabel space 4484 -3490 4484 -3490 7 sel24
rlabel space 4478 -2966 4478 -2966 1 sel25
rlabel space 4481 -2440 4481 -2440 1 sel26
rlabel space 4483 -1922 4483 -1922 1 sel27
rlabel space 4483 -1394 4483 -1394 1 sel28
rlabel space 4483 -877 4483 -877 1 sel29
rlabel space 4484 -351 4484 -351 7 sel30
rlabel space 4481 173 4481 173 1 sel31
rlabel metal2 3953 -17017 3953 -17017 1 A0
rlabel metal2 3518 -17014 3518 -17014 1 A1
rlabel metal2 3095 -17013 3095 -17013 1 A2
rlabel metal2 2671 -17016 2671 -17016 1 A3
rlabel metal2 2252 -17014 2252 -17014 1 A4
<< end >>
