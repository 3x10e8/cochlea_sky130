magic
tech sky130A
timestamp 1639217340
<< nwell >>
rect -371 527 1084 544
rect -439 519 1084 527
rect -439 450 1091 519
rect -431 -56 1092 32
rect -441 -472 1098 -468
rect -441 -557 1104 -472
rect -431 -578 1103 -557
rect -442 -1117 1092 -1028
rect -322 -1582 1083 -1519
rect -322 -1611 1088 -1582
rect -321 -1669 1088 -1611
rect -318 -2117 1083 -2054
rect -321 -2204 1088 -2117
rect -318 -2659 1046 -2588
rect -319 -2746 1090 -2659
rect -319 -3165 982 -3093
rect -319 -3187 1096 -3165
rect -314 -3252 1096 -3187
rect -431 -3839 -337 -3687
rect -12 -3830 82 -3672
rect -436 -4085 -257 -3839
rect -431 -4231 -337 -4085
rect -12 -4086 163 -3830
rect 410 -3838 504 -3672
rect -12 -4216 82 -4086
rect 410 -4092 587 -3838
rect 410 -4216 504 -4092
<< pwell >>
rect -162 -843 -21 -737
rect -113 -2359 -4 -2284
rect -139 -3447 -47 -3353
<< psubdiff >>
rect -162 -771 -21 -737
rect -162 -817 -119 -771
rect -62 -817 -21 -771
rect -162 -843 -21 -817
rect -113 -2298 -4 -2284
rect -113 -2345 -92 -2298
rect -21 -2345 -4 -2298
rect -113 -2359 -4 -2345
rect -139 -3378 -47 -3353
rect -139 -3429 -121 -3378
rect -69 -3429 -47 -3378
rect -139 -3447 -47 -3429
<< nsubdiff >>
rect -169 507 -67 525
rect -169 484 -147 507
rect -88 484 -67 507
rect -169 469 -67 484
<< psubdiffcont >>
rect -119 -817 -62 -771
rect -92 -2345 -21 -2298
rect -121 -3429 -69 -3378
<< nsubdiffcont >>
rect -147 484 -88 507
<< locali >>
rect -169 507 -67 525
rect -169 484 -147 507
rect -88 484 -67 507
rect -169 469 -67 484
rect -162 -771 -21 -737
rect -162 -817 -119 -771
rect -62 -817 -21 -771
rect -162 -843 -21 -817
rect -113 -2298 -4 -2284
rect -113 -2345 -92 -2298
rect -21 -2345 -4 -2298
rect -113 -2359 -4 -2345
rect -139 -3378 -47 -3353
rect -139 -3429 -121 -3378
rect -69 -3429 -47 -3378
rect -139 -3447 -47 -3429
<< viali >>
rect -129 489 -105 506
rect -524 149 -493 181
rect -531 -376 -503 -346
rect -107 -805 -81 -787
rect -528 -897 -495 -869
rect -528 -1414 -499 -1391
rect -528 -1940 -494 -1913
rect -79 -2337 -33 -2310
rect -526 -2466 -497 -2436
rect -519 -2980 -482 -2959
rect -113 -3423 -76 -3386
rect -514 -3512 -475 -3481
<< metal1 >>
rect -762 457 -556 761
rect -138 510 -110 511
rect -147 506 -88 510
rect -147 489 -129 506
rect -105 489 -88 506
rect -147 484 -88 489
rect -762 429 -483 457
rect -138 429 -110 484
rect -762 -66 -556 429
rect -533 181 -483 190
rect -533 149 -524 181
rect -493 149 -483 181
rect -533 140 -483 149
rect -762 -94 -477 -66
rect -145 -94 -117 1
rect -762 -589 -556 -94
rect -540 -346 -491 -334
rect -540 -376 -531 -346
rect -503 -376 -491 -346
rect -540 -383 -491 -376
rect -762 -617 -481 -589
rect -132 -617 -104 -504
rect -762 -1112 -556 -617
rect -119 -782 -62 -771
rect -119 -808 -111 -782
rect -75 -808 -62 -782
rect -119 -817 -62 -808
rect -538 -869 -481 -855
rect -538 -897 -528 -869
rect -495 -897 -481 -869
rect -538 -908 -481 -897
rect -762 -1140 -486 -1112
rect -125 -1140 -97 -1040
rect -762 -1635 -556 -1140
rect -537 -1383 -486 -1378
rect -537 -1414 -528 -1383
rect -497 -1414 -486 -1383
rect -537 -1423 -486 -1414
rect -762 -1663 -481 -1635
rect -53 -1663 -25 -1570
rect -762 -2158 -556 -1663
rect -537 -1913 -479 -1901
rect -537 -1940 -528 -1913
rect -494 -1940 -479 -1913
rect -537 -1950 -479 -1940
rect -762 -2186 -486 -2158
rect -49 -2186 -21 -2089
rect -762 -2681 -556 -2186
rect -92 -2310 -21 -2298
rect -92 -2337 -79 -2310
rect -33 -2337 -21 -2310
rect -92 -2345 -21 -2337
rect -535 -2436 -484 -2427
rect -535 -2466 -526 -2436
rect -497 -2466 -484 -2436
rect -535 -2475 -484 -2466
rect -762 -2709 -486 -2681
rect -95 -2709 -67 -2598
rect -762 -3204 -556 -2709
rect -531 -2952 -467 -2943
rect -531 -2982 -519 -2952
rect -482 -2982 -467 -2952
rect -531 -2999 -467 -2982
rect -762 -3232 -477 -3204
rect -98 -3232 -70 -3133
rect -762 -3860 -556 -3232
rect -121 -3386 -69 -3378
rect -121 -3423 -113 -3386
rect -76 -3423 -69 -3386
rect -121 -3429 -69 -3423
rect -528 -3481 -463 -3467
rect -528 -3512 -514 -3481
rect -475 -3512 -463 -3481
rect -528 -3520 -463 -3512
rect 148 -3603 229 -3596
rect -276 -3618 -202 -3614
rect -276 -3659 -272 -3618
rect -209 -3659 -202 -3618
rect -276 -3666 -202 -3659
rect 148 -3655 155 -3603
rect 222 -3655 229 -3603
rect 148 -3666 229 -3655
rect 571 -3610 649 -3603
rect 571 -3659 579 -3610
rect 642 -3659 649 -3610
rect 571 -3666 649 -3659
rect -762 -3888 -381 -3860
rect -762 -3975 -556 -3888
rect 129 -3863 211 -3856
rect -73 -3899 44 -3871
rect -73 -3947 -45 -3899
rect 129 -3900 133 -3863
rect 207 -3900 211 -3863
rect 553 -3870 622 -3847
rect 129 -3908 211 -3900
rect 367 -3906 469 -3878
rect 553 -3904 556 -3870
rect 367 -3943 395 -3906
rect 553 -3916 622 -3904
rect -762 -4013 -410 -3975
rect -73 -3985 100 -3947
rect 367 -3981 534 -3943
rect -762 -4142 -556 -4013
rect -283 -4015 -202 -4008
rect -283 -4056 -276 -4015
rect -209 -4056 -202 -4015
rect -283 -4067 -202 -4056
rect -652 -4272 -624 -4142
rect -652 -4300 -381 -4272
rect -73 -4277 -45 -3985
rect 142 -4015 223 -4008
rect 142 -4056 149 -4015
rect 216 -4056 223 -4015
rect 142 -4060 223 -4056
rect 9 -4072 326 -4060
rect -449 -4346 -387 -4300
rect -73 -4305 41 -4277
rect 13 -4346 41 -4305
rect -449 -4348 41 -4346
rect 367 -4344 395 -3981
rect 567 -4008 638 -4004
rect 567 -4060 571 -4008
rect 631 -4060 638 -4008
rect 429 -4344 457 -4292
rect 367 -4348 457 -4344
rect -449 -4374 457 -4348
rect -4 -4376 457 -4374
<< via1 >>
rect -524 149 -493 181
rect -531 -376 -503 -346
rect -111 -787 -75 -782
rect -111 -805 -107 -787
rect -107 -805 -81 -787
rect -81 -805 -75 -787
rect -111 -808 -75 -805
rect -528 -897 -495 -869
rect -528 -1391 -497 -1383
rect -528 -1414 -499 -1391
rect -499 -1414 -497 -1391
rect -528 -1940 -494 -1913
rect -79 -2337 -33 -2310
rect -526 -2466 -497 -2436
rect -519 -2959 -482 -2952
rect -519 -2980 -482 -2959
rect -519 -2982 -482 -2980
rect -113 -3423 -76 -3386
rect -514 -3512 -475 -3481
rect -272 -3659 -209 -3618
rect 155 -3655 222 -3603
rect 579 -3659 642 -3610
rect -291 -3904 -220 -3859
rect 133 -3900 207 -3863
rect 556 -3904 631 -3870
rect -276 -4056 -209 -4015
rect 149 -4056 216 -4015
rect 571 -4060 631 -4008
<< metal2 >>
rect -533 181 -483 190
rect -533 149 -524 181
rect -493 149 -483 181
rect -533 140 -483 149
rect -540 -346 -491 -334
rect -540 -376 -531 -346
rect -503 -376 -491 -346
rect -540 -383 -491 -376
rect -119 -778 -62 -771
rect -119 -813 -114 -778
rect -70 -813 -62 -778
rect -119 -817 -62 -813
rect -538 -869 -481 -855
rect -538 -897 -528 -869
rect -495 -897 -481 -869
rect -538 -908 -481 -897
rect -537 -1383 -486 -1378
rect -537 -1414 -528 -1383
rect -497 -1414 -486 -1383
rect -537 -1423 -486 -1414
rect -537 -1912 -479 -1901
rect -537 -1940 -528 -1912
rect -494 -1940 -479 -1912
rect -537 -1950 -479 -1940
rect -92 -2309 -21 -2298
rect -92 -2337 -79 -2309
rect -33 -2337 -21 -2309
rect -92 -2345 -21 -2337
rect -535 -2436 -484 -2427
rect -535 -2466 -526 -2436
rect -497 -2466 -484 -2436
rect -535 -2475 -484 -2466
rect -531 -2952 -467 -2943
rect -531 -2982 -519 -2952
rect -482 -2982 -467 -2952
rect -531 -2999 -467 -2982
rect -121 -3386 -69 -3378
rect -121 -3423 -113 -3386
rect -76 -3423 -69 -3386
rect -121 -3429 -69 -3423
rect -528 -3481 -463 -3467
rect -528 -3512 -514 -3481
rect -475 -3512 -463 -3481
rect -528 -3520 -463 -3512
rect -526 -3627 -336 -3558
rect -60 -3562 82 -3549
rect -276 -3618 -202 -3614
rect -526 -3895 -427 -3627
rect -276 -3659 -272 -3618
rect -209 -3659 -202 -3618
rect -276 -3666 -202 -3659
rect -60 -3627 86 -3562
rect 371 -3567 513 -3566
rect 148 -3603 229 -3596
rect -295 -3859 -213 -3852
rect -295 -3895 -291 -3859
rect -526 -3904 -291 -3895
rect -220 -3874 -213 -3859
rect -220 -3904 -205 -3874
rect -526 -3968 -205 -3904
rect -60 -3899 30 -3627
rect 148 -3655 155 -3603
rect 222 -3655 229 -3603
rect 148 -3666 229 -3655
rect 354 -3631 513 -3567
rect 571 -3610 649 -3603
rect 129 -3863 211 -3856
rect 129 -3899 133 -3863
rect -60 -3900 133 -3899
rect 207 -3867 211 -3863
rect 207 -3899 218 -3867
rect 354 -3899 445 -3631
rect 571 -3659 579 -3610
rect 642 -3659 649 -3610
rect 571 -3666 649 -3659
rect 553 -3870 638 -3863
rect 553 -3899 556 -3870
rect 207 -3900 220 -3899
rect -60 -3968 220 -3900
rect 354 -3904 556 -3899
rect 631 -3882 638 -3870
rect 631 -3904 642 -3882
rect -287 -4008 -205 -3968
rect 136 -4008 218 -3968
rect 354 -3994 642 -3904
rect 354 -3998 445 -3994
rect 564 -4008 642 -3994
rect -287 -4015 -202 -4008
rect -287 -4026 -276 -4015
rect -283 -4056 -276 -4026
rect -209 -4056 -202 -4015
rect 136 -4015 223 -4008
rect 136 -4019 149 -4015
rect -283 -4067 -202 -4056
rect 142 -4056 149 -4019
rect 216 -4056 223 -4015
rect 142 -4067 223 -4056
rect 564 -4060 571 -4008
rect 631 -4060 642 -4008
rect 564 -4064 642 -4060
<< via2 >>
rect -524 149 -493 181
rect -531 -376 -503 -346
rect -114 -782 -70 -778
rect -114 -808 -111 -782
rect -111 -808 -75 -782
rect -75 -808 -70 -782
rect -114 -813 -70 -808
rect -528 -897 -495 -869
rect -528 -1414 -497 -1383
rect -528 -1913 -494 -1912
rect -528 -1940 -494 -1913
rect -79 -2310 -33 -2309
rect -79 -2337 -33 -2310
rect -526 -2466 -497 -2436
rect -519 -2982 -482 -2952
rect -113 -3423 -76 -3386
rect -514 -3512 -475 -3481
<< metal3 >>
rect -1179 192 -835 748
rect -1179 181 834 192
rect -1179 149 -524 181
rect -493 149 834 181
rect -1179 142 834 149
rect -1179 -331 -835 142
rect -533 140 -483 142
rect -1179 -346 840 -331
rect -1179 -376 -531 -346
rect -503 -376 840 -346
rect -1179 -381 840 -376
rect -1179 -854 -835 -381
rect -540 -383 -491 -381
rect -119 -778 -62 -771
rect -119 -780 -114 -778
rect -126 -813 -114 -780
rect -70 -813 -62 -778
rect -126 -817 -62 -813
rect -126 -854 -76 -817
rect -1179 -869 831 -854
rect -1179 -897 -528 -869
rect -495 -897 831 -869
rect -1179 -904 831 -897
rect -1179 -1377 -835 -904
rect -538 -908 -481 -904
rect -1179 -1383 842 -1377
rect -1179 -1414 -528 -1383
rect -497 -1414 842 -1383
rect -1179 -1427 842 -1414
rect -1179 -1900 -835 -1427
rect -1179 -1912 829 -1900
rect -1179 -1940 -528 -1912
rect -494 -1940 829 -1912
rect -1179 -1950 829 -1940
rect -1179 -2423 -835 -1950
rect -92 -2309 -21 -2298
rect -92 -2337 -79 -2309
rect -33 -2337 -21 -2309
rect -92 -2345 -21 -2337
rect -92 -2346 -22 -2345
rect -86 -2423 -36 -2346
rect -1179 -2436 823 -2423
rect -1179 -2466 -526 -2436
rect -497 -2466 823 -2436
rect -1179 -2473 823 -2466
rect -1179 -2946 -835 -2473
rect -535 -2475 -484 -2473
rect -531 -2946 -467 -2943
rect -1179 -2952 831 -2946
rect -1179 -2982 -519 -2952
rect -482 -2982 831 -2952
rect -1179 -2996 831 -2982
rect -1179 -3469 -835 -2996
rect -531 -2999 -467 -2996
rect -121 -3386 -69 -3378
rect -121 -3423 -113 -3386
rect -76 -3423 -69 -3386
rect -121 -3429 -69 -3423
rect -528 -3469 -463 -3467
rect -120 -3469 -70 -3429
rect -1179 -3481 853 -3469
rect -1179 -3512 -514 -3481
rect -475 -3512 853 -3481
rect -1179 -3519 853 -3512
rect -1179 -3847 -835 -3519
rect -528 -3520 -463 -3519
rect -1179 -3934 793 -3847
rect -1179 -4150 -835 -3934
rect -913 -4266 -850 -4150
rect -913 -4321 757 -4266
rect -913 -4349 -850 -4321
use pbulk  pbulk_7
timestamp 1639210801
transform 1 0 -438 0 1 -4014
box -18 -18 119 75
use inv_customized_3  inv_customized_3_3
timestamp 1639205400
transform 0 -1 45 1 0 -4223
box -85 128 180 481
use inv_customized_3  inv_customized_3_0
timestamp 1639205400
transform 0 -1 45 1 0 -3823
box -85 128 180 481
use pbulk  pbulk_8
timestamp 1639210801
transform 1 0 6 0 1 -3995
box -18 -18 119 75
use inv_customized_3  inv_customized_3_5
timestamp 1639205400
transform 0 -1 468 1 0 -4224
box -85 128 180 481
use inv_customized_3  inv_customized_3_1
timestamp 1639205400
transform 0 -1 470 1 0 -3823
box -85 128 180 481
use pbulk  pbulk_9
timestamp 1639210801
transform 1 0 431 0 1 -3988
box -18 -18 119 75
use inv_customized_3  inv_customized_3_4
timestamp 1639205400
transform 0 -1 889 1 0 -4228
box -85 128 180 481
use inv_customized_3  inv_customized_3_2
timestamp 1639205400
transform 0 -1 895 1 0 -3823
box -85 128 180 481
use 0  0_23
timestamp 1639200303
transform -1 0 -178 0 1 -3658
box -89 43 336 566
use 0  0_18
timestamp 1639200303
transform 1 0 0 0 1 -3658
box -89 43 336 566
use 0  0_19
timestamp 1639200303
transform 1 0 425 0 1 -3658
box -89 43 336 566
use inv_customized  inv_customized_7
timestamp 1639201766
transform 1 0 951 0 1 -3661
box -194 128 180 481
use pbulk  pbulk_6
timestamp 1639210801
transform 1 0 -129 0 1 -3172
box -18 -18 119 75
use 0  0_22
timestamp 1639200303
transform -1 0 -178 0 1 -3135
box -89 43 336 566
use 0  0_16
timestamp 1639200303
transform 1 0 0 0 1 -3135
box -89 43 336 566
use 0  0_17
timestamp 1639200303
transform -1 0 672 0 1 -3135
box -89 43 336 566
use inv_customized  inv_customized_6
timestamp 1639201766
transform 1 0 951 0 1 -3138
box -194 128 180 481
use pbulk  pbulk_5
timestamp 1639210801
transform 1 0 -124 0 1 -2637
box -18 -18 119 75
use 0  0_21
timestamp 1639200303
transform -1 0 -178 0 1 -2612
box -89 43 336 566
use 0  0_15
timestamp 1639200303
transform -1 0 247 0 1 -2612
box -89 43 336 566
use 0  0_14
timestamp 1639200303
transform -1 0 672 0 1 -2612
box -89 43 336 566
use inv_customized  inv_customized_5
timestamp 1639201766
transform 1 0 951 0 1 -2615
box -194 128 180 481
use pbulk  pbulk_4
timestamp 1639210801
transform 1 0 -73 0 1 -2129
box -18 -18 119 75
use 0  0_20
timestamp 1639200303
transform -1 0 -178 0 1 -2089
box -89 43 336 566
use 0  0_12
timestamp 1639200303
transform -1 0 247 0 1 -2089
box -89 43 336 566
use 0  0_13
timestamp 1639200303
transform 1 0 425 0 1 -2089
box -89 43 336 566
use inv_customized  inv_customized_4
timestamp 1639201766
transform 1 0 951 0 1 -2092
box -194 128 180 481
use pbulk  pbulk_3
timestamp 1639210801
transform 1 0 -82 0 1 -1610
box -18 -18 119 75
use 0  0_11
timestamp 1639200303
transform 1 0 -425 0 1 -1566
box -89 43 336 566
use 0  0_2
timestamp 1639200303
transform -1 0 247 0 1 -1566
box -89 43 336 566
use 0  0_7
timestamp 1639200303
transform 1 0 425 0 1 -1566
box -89 43 336 566
use inv_customized  inv_customized_3
timestamp 1639201766
transform 1 0 951 0 1 -1569
box -194 128 180 481
use pbulk  pbulk_2
timestamp 1639210801
transform 1 0 -153 0 1 -1085
box -18 -18 119 75
use 0  0_10
timestamp 1639200303
transform 1 0 -425 0 1 -1043
box -89 43 336 566
use 0  0_4
timestamp 1639200303
transform -1 0 247 0 1 -1043
box -89 43 336 566
use 0  0_6
timestamp 1639200303
transform -1 0 672 0 1 -1043
box -89 43 336 566
use inv_customized  inv_customized_2
timestamp 1639201766
transform 1 0 951 0 1 -1046
box -194 128 180 481
use pbulk  pbulk_1
timestamp 1639210801
transform 1 0 -164 0 1 -545
box -18 -18 119 75
use 0  0_9
timestamp 1639200303
transform 1 0 -425 0 1 -520
box -89 43 336 566
use 0  0_3
timestamp 1639200303
transform 1 0 0 0 1 -520
box -89 43 336 566
use 0  0_5
timestamp 1639200303
transform -1 0 672 0 1 -520
box -89 43 336 566
use inv_customized  inv_customized_1
timestamp 1639201766
transform 1 0 951 0 1 -523
box -194 128 180 481
use pbulk  pbulk_0
timestamp 1639210801
transform 1 0 -177 0 1 -36
box -18 -18 119 75
use 0  0_8
timestamp 1639200303
transform 1 0 -425 0 1 3
box -89 43 336 566
use 0  0_0
timestamp 1639200303
transform 1 0 0 0 1 3
box -89 43 336 566
use 0  0_1
timestamp 1639200303
transform 1 0 425 0 1 3
box -89 43 336 566
use inv_customized  inv_customized_0
timestamp 1639201766
transform 1 0 951 0 1 0
box -194 128 180 481
<< labels >>
rlabel via1 181 -4044 181 -4044 1 OUT
port 1 e
rlabel metal3 -1016 731 -1016 731 1 GND
rlabel metal1 -659 739 -659 739 1 VDD
rlabel space -255 -4258 -255 -4258 1 A2
rlabel space 173 -4257 173 -4257 1 A1
rlabel space 592 -4260 592 -4260 1 A0
rlabel space 1122 281 1122 281 1 Sel7
rlabel space 1124 -238 1124 -238 1 Sel6
rlabel space 1127 -761 1127 -761 7 Sel5
rlabel space 1127 -1288 1127 -1288 7 Sel4
rlabel space 1126 -1810 1126 -1810 7 Sel3
rlabel space 1127 -2334 1127 -2334 7 Sel2
rlabel space 1127 -2857 1127 -2857 7 Sel1
rlabel space 1127 -3380 1127 -3380 7 Sel0
<< end >>
