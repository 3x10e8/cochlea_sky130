magic
tech sky130A
timestamp 1639210801
<< nwell >>
rect -18 -18 119 75
<< nsubdiff >>
rect 0 45 101 57
rect 0 14 21 45
rect 82 14 101 45
rect 0 0 101 14
<< nsubdiffcont >>
rect 21 14 82 45
<< locali >>
rect 0 45 101 57
rect 0 14 21 45
rect 82 14 101 45
rect 0 0 101 14
<< viali >>
rect 36 21 66 38
<< metal1 >>
rect 21 38 82 45
rect 21 21 36 38
rect 66 21 82 38
rect 21 14 82 21
<< labels >>
rlabel viali 60 29 60 29 1 Out
port 1 n
<< end >>
