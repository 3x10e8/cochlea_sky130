magic
tech sky130A
timestamp 1639201766
use 0  0_7
timestamp 1639200303
transform 1 0 425 0 1 -1566
box -89 43 336 566
use 0  0_6
timestamp 1639200303
transform -1 0 672 0 1 -1043
box -89 43 336 566
use 0  0_5
timestamp 1639200303
transform -1 0 672 0 1 -520
box -89 43 336 566
use 0  0_2
timestamp 1639200303
transform -1 0 247 0 1 -1566
box -89 43 336 566
use 0  0_4
timestamp 1639200303
transform -1 0 247 0 1 -1043
box -89 43 336 566
use 0  0_3
timestamp 1639200303
transform 1 0 0 0 1 -520
box -89 43 336 566
use 0  0_1
timestamp 1639200303
transform 1 0 425 0 1 3
box -89 43 336 566
use 0  0_0
timestamp 1639200303
transform 1 0 0 0 1 3
box -89 43 336 566
<< end >>
